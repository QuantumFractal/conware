XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P��:��u��)�$l˾�=��Y��g`D��ۣ}8}aoN^J�y���"�𔽖�������lk����tl�;
���ɵ�V���v�%��4ɷ��iv�����UI9�>CQg��?�SZ���~?v3�#�E;}�w�ID�S�4#Q[u��y3v.#~b�X���y���3�Ex�d�.	Yx��;.�\V�����$��U���{�Pw�������)��2K���cb�@i���~6�*S/~��0Ѿ��-f˱�J�̿���C�'X�p�Ӆ(::a�6��c�z|�M�p¹���$K=�>��k+��֧-��T`$�b~ݝ�[�S�N0!d���7���B �_1lU ~:��O$�J�˿��ǚc�hV/�
qo���J���ˏP<f��`�<�:f_�#�X����%Ϙ�XxBU;9�I�Փov��[\,��K���IL�F�MCp�N�d��W#�� aY$1�����U��͎b�t�/���TȨ2��ذ0 �RY�s���b�Z8��S�4�Z^��N4��o�!y}q�(<����a���n�H�~U)�p�̝L�C8���em����v4LK�H��^�6׫n"�<l�g.�E�<_��o7R/up�:�:��0tS���˫��?�{�E��� I{VZ0����1L!�X*x�8(_�o�"( A+H������fZ�:/���CZ(�I��ۘ�}�ϣ���ce�s�m�F /p��#H�,�/q�t9v���jѝ��Q�d��A��XlxVHYEB    b3c6    25b0h�"�u*4?���!
@v,�DDCG��0�ڢ6���Y�JHI#�6�_N�
���}��*�P:��N�?��_E�������T���E��p�:ت������Gn�M���<��;9;�%���ݯ9R���&��Ԁ5�P���(Il�sa�8YSް`��C�u=1��h��͑��5k�/�?�(@_�b�� �^V��4>(?k���)��Z^�i��Uxa6�|N.�R|���i��MS3�u��;��igfc)��vFg��k��-.!ló���~�{�*Cb��}�
�����NŽ?4�\A2� C���� 5l�RRtfӁ�V��㸺:��_*x�u�eA��_@	51Zq)�j�?������4�v��$Jy���_U탨j��:�ASB���4�M�TH5)g�he�&C�-H=���H���y(n.������#oǦ��J�����By �/6a��P�ˡ���x��&>�ȣ�oe���Ӆ��+!�jb�c�1uN�?ƳV��m���\����U�/��M��H�^�vZ�ލcw�%��i-r����`z|pS����č��1`�]A��s�>��TlI
"	!��q6)I�Y߼{��ʘr��v?C��)|��D
Xa�N�OM�L��<
C��E�4�
C� �Z_�u� =�Ai����$�"���N��E&i>N:��M�>�!m���ASo3��E��9���� �*M�V���ǻ]��C7��lX[k��o��� ^ZSg���߄����6!6N�"���gH�R�9K�ybo�) ��Ơ�}��ʨ�%�.�a?�gD����Un�HGF]#7���Gx�R^j��������Hn�~����8���D�
IL2N��8C���*\�^Gc�-�Dp���{a"��QyQ��u�x>W�;LQ���7X�ߋLOc�t8��w*ڰ� ��ۿ96D鋇�Z?OGo@*)�씡t`.�(b���q�R��#�a�z�p�uR��$�3�gS�9^RW���ǒ��-����|��ʨ�<\p�/�_�c�f���.{��d���A���,�,`pXf%߼��pt]j/`��J�a�L/++����������=s7D�����u	zd�az��mW�2z�|`s�����`5�:��������wkMP=f(@�㶎{sw<�q��W���?���#��橚&���O}>e�)_�`[�I���A�ѕ��a�q��7�����m��J�RSJ���z��Ra�σ��y�x�������Q]}W�'%��y�����~���"�K���<i	��K�4/L�=�9Ȏ���;o�A������h�?���p2�%�>��VҔ�t:�q�����x�shtyRWW&|@l��:"�,M����S%��]-� D��Lƥ��`^��E�%�*���)l��	U��u��IB��do�l���F�cxͤ���'V���8\�pk�6��F|�Đ�C_p%)|\�'Uc���Zx���L��j[p(�t� �N�q���~�Iԍ	��Ay�,��;�Aw	���+h:��j�a�NV!D?�˷.M���,Dn�ٚEj&V�aQ��$��	F�����O,��Lj�{E�W�����ESZ�G�zŽ�޵K`TuVZs���Z_�g�1�i�]�%&�mnܱ��1�,CKGYn|�䉒�bNg\�;��n:�O����A�c�m�����z��<Lf�*�D���&< y�0sH��h�^�l�F���F�����[���p�ߺu"|K<��F?V�g�'f����ډKy|��މ�EwiP��Z���#��e�<,�p,i�������lb��,X�R�7O�]I�&�?OP�>�aJE~&:6k�_,�rc}�xz�1ʹ�]�ղȟX3R��
�78&��U���!�k�ҽ��c��zb�m��&9PG��ȉ�F��u^�F.�|@Klm?�/��e�0v��%�(I O�;鎃��,0SOcF���<����Q����՗Ǘ+ۘ�9����@H8��D���BR�7�� ���B���J8pY�G@��ƞ���34�0^eW.���/nos�LU�%:���X8��`� I�<M�؝�����Y�+ �E��E��U���q̵��%��;W�F�M[y�f��$�Eg�Kz;>J�Z�ƏN=r��r �4޾81�?�)-���;8W�2�`ƻ�=���Z1��M�p\������
�]l�ꫮ����g��6?�����&q?�87�������l3q��ͤ�Ǝ�,�h�U��wz�,h�`����{��t���ɔ"Ò�p��TUAԁf��0�u�EȚ~VǢ��6�o wY��iA�8��a�Ϸ�����'G-�Gt[�E>���H�����{4g$�-�v
٠R�Ɏ[��
�dz�h;N��:���Ņ��j��4?_���8�}�V�v���U�<'L�G$�#�c�����hd>+9�� ��[��	` �y�5^�*	��Z�)���B�=#B13Z ����Ш��v�b�t���}R����v��
�#�H��[r����{u�j"�j�h.�ʞ�3�$���l?Z=��B��sÐ��qOv)�����a�s|��n�{�u�[��]���3�=W�z�#�PY?Ftq��b��/���,2���S�G9�����Ņ���6�B�n�R��IU��L�M·/�*�{Oͬ�p��ɶL�����A�|���P^w��'�(� 
�R�
S����y�0���bw]�>)4e�:���_�ԟ�Y�Ȯ|0U(��A�m��c�T�6�zɱn������⒠f[y�#�-*�9�Tn|��d�T7xg�2�3����8��˫xi	7
����JK��-�����%lI�-���&Uk��8��䡹�J�+,�C�;��~M��Q|ڔIDM�������'��Ez�R�ob���3o�.�,�*nK!8�[~��v=)9�8�=�%��S�P���*x>�Ò411dIV�������<�j�Id�����X�h����3U�p����=�.������Sdj��z:��)o�>��H/�Afӱb&����/�G��!�=�w/k�w���H��dj�C	n�Y<k�L��l����a��?h�T@݌�J�
��n+�ޭ�MJ�#����&дn��(��6��X'`k���]ߵ�(�e�lP�e���A/��	6fX_c>9����MB��B�t5��е���ф.0S�|�4T|(�"�UO߱�7��&�,�����\�KQ'�m-����Cy��B'�c�Z4P�>Ļ��?���4uR<u�\n�_�5*�!c��m����:�����S�����7�y&/~YD�wRG��#,�PHK���X4x��ey��Ӂ�&;M3�H��I�q��Dn���hS�Y�.�1�噷vx��� ���d�����v �,�^��� ���H_7�7'�LٜW�`�uDӱ*]w�\��m�<?��jo���續/�o�� `<_��F��|��gY�O���$���9Ο��kjZ��:�GC
�"�4����T������pX]vh�N��&Z���p�������MN�9�1ь�/Y�߈��6��V@���K��T�����V��S�*�ŊT�@>O�
km�!��E��pج#R���F�byS��@� �0�"�B�I-�*�ڊKl�ٌ�vv��������sÙ�[M6�� ��WΈb�i:���S�mPa�4�W`� � ֮�e�����)W :RMG�e=�L�ST�WУd�Z�2a2�B��Ukg�e0�;|y~�ba����a�����Y��]6a W��5�b$�}�կ�R�8�RK��V��\�a�~�`Mi,���9��ŶV���B��ef��ko(]�D`t{��������J{K�4~.T��(��-qa��\�m��w����R��*j��c[����#8J�u��M�ϟ�ǐ#�P���Z���Q�����9�d뺴�� �������,/A���dh����r��DlP�]��R^�e�S �shZ8n���g���5���E��k��Ęh=��L=V@<' \�|�c�lC�t}���t�t�+���K�eU)�eH�!=%��؉H��~q�,@����+磺�^`��{l�ni�������p�����P�_P6��Xː�s���
e�H+�dˋ�r#!$��|��_j#��l�$x��"�����b�!��i�M�$Эju�{nuA�P\.x1�+:�`�s��	By�)�/�[=�Z���������ښZ�P�0����b���5R.gv:�F�ٺ�oU���/o��Ψ{E��H����U${׺�y��uNҲ�rԘ7�
,��H:���g�����v:�ohAJ�g7�X�i��������e8ˌ')s��-�b�e5ĝ
�6}}�T����[��u��s�d{_�����>S�����Z+��5Sе��	�����Wޅmj*�K.��i��@�ӕV�櫓�Y�~d���3�x���f�����΋ �Bi�2�~d�Fo� ��H�6r�s!����&��5a��q��k�F���%r��:2Q���W[�7��>۶`|��'ع�� ��(���� ���p!�s�nǤdr���UC�����"
���9��l��k��Y�eO(����M���e��<�&AL�Wr�tJbmR���������)��q�.1@����筌�p�x�u�G�"���x��j�Ek���3���MP���Vv�M�e����4�d�>bDANj�.{�eUC�o����9~Iq��z �#w&P=�)�M��5p��;fmz)���q-����[KB �n��)���������"���Y�-��h�{Iu���?%4{�����a+t��&�s��$пWutCD:��� H�E�xB��'K�O(l��4GK�Ć^����J�z$f����,�<��2$��|���R1�j�	��J��PU1�J��''
�� �W!+</�B�j�+c��ʺxO��Z	���M�0�Z���ǧ�^���}�*2}�9 ����u܏��%��ZZ=��L#�L�J�՘�&���4X��.�l('B���i<��!��$�ƹ�����1�P��Lwٛ�#� V�Ļ�A�h,=��P�P�y|�#Q9٧$�fB��A��vl�=���DXS��0���7.����
����!:�nZ���
�r�Q��8��TȨXF�6�3{�&��7O6�y��2���։*�����*���/RX}F{uy_�dE��+��^�誤���'�קƠ�KLR�hiԷ9�=Y�����po�dQ�J�0,�%^;������7������m��-�4�8*�������Y�WL*qh<1��)�Hc|�߆m�}*Ye�G-�k.����O�	w_��V���Ì������(����|�{Q�
�Wʵ�7}�?)р�I�L/$Io��H�9�HC�Vo��O'S�}����C'�g�S�P�.0ԯ���%Bם`='��`n�7;x��h�H�N��T��1��NƎ���<����">v�7}�`6�e"ɕ��/�:�-H���\�h"p%����3��f?�Q����"�F����Y�ڒRs�sx�LoY��,�����M9m��C�@��a��P˵_G�arN(�Y<�NH"hVix��UF�o���Xr�:��Ozz ��ݞ�zu��XUK�'���<�f�Q/8�&�ǏA��)0�TTTq�PL�╀-$`��YP���{��v�p�)���j�L�6B��L^5h��c���d;�4#�1<�.V{�ɂ���1N�YN\�gv���Ѳ�/��P�@Ɂ����ՙ'�67���z�r�}ߎNG�0p�ԫlR�$w�L~		V�PĪ!��S϶���%*��m�~�NI���9���%n}�M�W;�f�ߠ�Xk�K��ޙ�Q�b�(4l&�;=�����J��x%�
/��ùհ�j����Q󉊹6E%-����?B�7+*&���1E$%F>�c"9JoBa��C1��Ao�!�&>7��rU��.�Tu Y&
Qzd���/6v��y�7��"���.{��*<����*�/���e��0��s�����qnp�� �R���KpȊ����bz ��[!����X��_��mw���"Q�~��)d���rd�.@a�+'�􄐁��s;��'ľ�#�:dǑ�a�أ7#&��6js7���nߡ���ϒ:&Ϣ4�|�����y�HB��*�e[j��/f��-�J��]5�=��7T�b+Y�`.����ޡ��'���2��'Cg��0Q��J1��(�03�G��ǩf�i,��ej::��fRR"7:�o?3�(�r�yD�w0F�R}�I|�O��ӵ�^1���0�o�#W!� �+�
,A�jV9�D��ı3)y��K�?*�{?A�Y%[��k϶[�����R*��΃�.��s�h��k,�_f�BJ�BA(����:;�ΉZ�W����lU�C�F�B+-l�]�&TLN�HɵA��{f�9-C4h�![�qY����/�G�h]����g��_�Ř"�%9�u��m��[�,�y�,��>=T�`?DhyZ�mۓ��$R������Y���Ji�A)(|����}�#X\HC	0[�!�8�E2?!�	&�߫~�j&�1��� �3��<�{�6�i�]]����Y(|ï�'�pJiT�7�)�^1�>�u�o�.�׷�ۻ�b�[A;���Dv/�S��'���,Z�7�@����4x�>�%$�X�)a�dY���0-���r�=,��G��2|��AD�����'N���h��M@zpk���!��b���_�6�8(_��d�ʏP@Z��Co�F�$g%���w���,��J�B��4�&NC�e��+�R��7P���?A�z��u�*ߊ1��z��ڴ����-�� 7Q�&b2����j|����q%CX��>Y57�,�8��v��[����� �`����FD�O�I�6��EoC��^�e:O�ۆ�M �|c�ׅ��`X���Y��s��4��@[������=��0\;�r��a�D�ⷭ���Á!��_J�����e�M�����)�3��3@]�bO���" Y����"=� q�4��`E����
0=	KDV����ll�mB덵~J%��MRy������Πf�*	�6/�BP}�RF|:�+i��ċ�]��228�"j�jW�Q;�$���M����x�#�[r�"B4���%cR�ҹ�ܗ�n���m�#��Nͥ���^�s���׺��5W�����ޏ�u�Eqy���7�tܐ$����LF��uY�6}gG�G�ob_��祬�TJj]�F�Rȹ�D�֨�T�D���U �cN&�?���.����2��	�Ll�{�c!�7���Z��fb�J96WE��m]Ё5bLP�6�����,��5�+��6�hK�fdX�j#�|��nW;t31��'2�
���%]�_�K�y`5���k<m�%풷Ҫ�5a���'��,#/��)V� ]�Q2����nJ��!|l�ʇ�f��E���jI��V�TKl���;�},}����s@6���[��R�圩�M��L8��F(�ݓ:I�S�����/(�N��Q�ĕi�ߜt�-���/x�xu�P5̄8�������(�c[7�H*��tsI7@?n�	�� �c:�>��Wfr��\3Թ��wd<�o��9��sj7�kò�����>l�x�M���.~���0$�7t��bP6�M�����vV�t:��%u@u��۲c�V�H9�O�*x�n��Li�eP�����C`�4�Q�Ĩ���rJӄi�p�C< 'Qq4���̫W\W��*|��E�˄����A`�ɇ^��P'7.f�������Ûvv����{FG�n�����������\ )|��p�е��3��" K!��e�F�0�����6�n^��	Yb�󜕸^�!�����w��G�����+3,7.�f�b�$�Q�^>��/�<hK^�A�ğ��:��Z���%�;U�wK�D�`��e����C%�{ٶ���e��@������r�.l��Y�3�f�����}�@L>;^c�G�뻸6v����Ն������ع%$�
-�o��� ���pO[� Vs�pC�}�Bi׸�M��f���;�?#7���6B���x!��9������V�Y��'�M&�M��t^�9ꢒ���;��ȗ<u�����r����Ph1�I�(�?Mc��K���TcS�{�N�����a?�&ȶz�F�PpY}��r�u�?��Ct�C:T��fF�0�g:Cb���"hON�X.��٘hT5����n����t�n+4�B7¹��5(�Ô4�̶��p>�0*�)k�saS�RR��Wv���5��ԅC�j\MO�J?k����T=�jqW�Ow�>"*�����	-	m)���W����F>q�x�Q�zϝHgt��i��;���&V� H�]�����l�t��d��+1��5�x��C˴���U��*��� ���v�Zy_T���#��#�[��x�+:M0jt쉮����ʣ#�*e�U��+/çL�'�
���_S>o��fi����\\�['�^����B�\Y�Y��z�3&���3���tT�L����M�QR��+���pJ��������
k�݉]��g��1KLeqx�U��g;B0DnA���*���`��ן�a��n�-�������>�3%�хO��T�\"%�sR�����ԓz�\s��/�!���M5%���8���m�+uf�OMY�W�ؾ��oa�r���In��"c��=/��m%���]`Ր�R�E��dל�RG��cM�j8�����
HYZw��$a$�Z�\�U��mȈ ��ח%!�������~��GJ�l���ISJI�*p����U����i^$-�h$(���v,}<�>.���*�%��M��"�Ť��艘V�{��x��+���7�0��8�-=a�i-E�2���#��KRA��UF�]�]��u��)���Yjʅ�f�bj�Т<I ϴM�8��Q���]����G�֦�
!�>��i[nu��� �0{թ��!�?�x��ڗ�

��n���ޞV۩,��ʺ������ҡ�\�5���XJ!��j���Ҏ?��ǲ ,r�㾗f�8��4����s�s��[\�Ne���r+��n�^�ti�Au�x���C��7^ ܜ�3�͖"P���d2����2�R�ٯyz�*7��"�:���p��	GHc7x@��~[���A��bӃ�o��X	�I�&�̴�>�ԧ`��)����Y��e�wo���Gt��{��>�a;&�KD�*�+�tCߖ�{��uK��[���]�u)n�3R�5Ix~��Nu�Or��l�ټB�� ���:�����nns{��U8X�hM���k`~}�mu������'�4LC��S�b'�
�#�N\<L�iq�l�4����8R�T�sg���'�/�sQS��