XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����Z�4_ѫ�<'�O�S.Xj��0���р����%�g�o�K-<2L����. �-��IIC��e׳̣돥g�����M1��φ{'|EC�̴�����Ȝ4$��g!� �.�����u.�b �L(�z�����f��H���	m�pl)ɴn|'��F��}�YpG���&47�.��-�;��l(oX��9�'�B�����	����8����Os:/�8]s�šd�G%��$�����~�u�:x��5���(��"y��h����42��!�#��y�1S�ο�_PG��.Ӳ�P�F�jZ�i���F���߻��GoV�ߑ.5�o��h.pF�R'�SL�Z~�o[#��V���\+y���@�惫��hRq�`�:jhw��!3g���=�9o�q�,)�A�~�So��=�㔠'4���&w�&���{����F�y*pzIO�4��9\��t3��D���zf���hB�9�m%�4�]�M�jX��P�ˆw1���nҤ�_��,���p�g?Z7&Z���[���\N�lȞ��RYw���R�L��妏�9JA���;n��S�av�-��e�d�^3 =�	��n��1U��E�P�Uy�#n���.y��3�D�3�����ԘWMD�ۿ�mɢ{��n~��Î��Fc��OY6�V ��n�p$���toP8:�ٍ�ΎS��uI�5�������i�f��|{S����5��7���%}ъ9��Q�L�x۲�Մ\�Ƽ~ʼ�֚���O�>��^i�p�ՃXlxVHYEB    dd8f    2160����.��yW�#�TTU��E$��+\nT�_%|��g����W��>�y�ĀUT��v|�4~�V�R^�����b;]��U��)�ѹ��O��D�$���3��VEu/,��
l���(y��Y���	����o2ɄΪ��8���Eiͼ�F�"l�k�\d�j�>rZv~�:A��p$ͯ{��gc�dG������w�
�մ>F�ι�sj����Ľ��CҺk�gB'��c�Ĺ�X\t��2	�D�&�ʚ�Yn_�B-�#G���{��P�� Tp�w,R�l���U҈�Cq>���e�oV�ձ�'w����v�����t!�{�&�,P�.�Ffa|)mD;5t֓3��R�!��,���>/ ��B�T!w7{�bJ�L~	+םp\����Z�+����I`Q���[�2�D�9}�ש����՛�T%n�Z�s��i_�[H;B�4���4�Y��OB�˾̾�6W��EPc��Q��E�N�$�\8g$ٺ�{v�K��9�"����B�Q�x��F���P6���56x�zo�v�WC�CU�k��h�U
=!���V6�"ެ�?B�%,��9/חG9A�	��"����^ş<!�<䝣��9��I r�=iJ�C'u�i��]Қ��Q���X��H��ҽ�Hk�����n~��fT�d��Vs}�H�o5����d}e�Hv�i5E�p>�CoF�*�V�W|gݳėJ1�H��A�����<��)6X�y&���X}S7�����p��r6Ü���g�'e$�Ox���bH��u�Ü���[�aW�$@� �r��,^|c(r�g|��#B�2���w��Ӑ��{P��BtC��_�I�iYf̜+�,��7�d�S е/�G�5q;Pi�˰颶B����-&���d�A�D��� �8�䬍z�׉!sn����΃1o���E�1l�O9����
l�s+�9���p�����/6"�����Z� k${M���(�ä�DL���i��[}���	;�%{��G4�t�m��2���b���>��豏g�ۺ��ۓ�R�����CP�ʲ���Pm�s֧8i���b�����j�X��YX���)ƞ�_C��v�+�$�i�_I��o��.��Щ��������]��^���j�4}t��q0V��+�]�-����I�+ϗX1���[T?2�n��آ\�:g~,��c�s;/0-�$��݂�H���!h��\����x.Ά@/a�r@
:E��JG�$��;Ƿ�g�����3�r�@")��K��|B�w�9v<��ŅJ�zQ]g|���V \���#�������r��ۡ��U��2+�G����HE��4�\�>Z|�u���.A�z'��O�մ�\^+G�~<��(%{��їSBaҔH
��>��g�(#q�ey&^+��u�r�c��iZ��²��fx��5�t42X�Q�
u��`�5ez���y������<��_�����Y�ӭ�q�����,�'�^37wh��-8��/u_ ҥ�3j:�?�,1z|0��G�5�=f�dI�w��@4�&��v���?�O���h ��5�Þ >f,C�~O����g��֭P�n\1r��V����:$�y�R����1М���f1}�
�4�,���,p3��/�=�Peqܣ��֎�XZ
"Rŗ�[��qrg�r���5Gw"A���,=��5����`r��n�Y���_ג7�ti�����hiͨ͟�&�4X�DO��NR]6Rt�Ĥe1I� ��m��Yy�X�}&o�6MWI�J�j����K���A�I3�VmNo��|{�j��ss&<4�fj�[�R�q#��cy�E�b�{����� �5�a{q����/5f�\�!TM����.��*�<S�Z�������i���s���]�QA�`(��/=�WS�E�ޣ�_�����j{���z^�@$ �r*|���0w�����1f�c�����7�����;[�E��7�i�K���/KǱ6(ܜ0͐���甁8%;_$����7ަ�L���@h)~3����%�x�-��~h}��l��L��#� ��	jQ d�^�}�C��ޕ�"�b,p#ei�H𼧭�C��j{D-N�:�FO��'��b.�#N2a�ԏ�|�z�v 6*���b�ٽt82�>[@��׍����.y��-���-�w��Z��v���z�p����#w�K���ɛf�y[oƛ.������s
�W������6�}�]��B�c������5 )H��RmHț����5����Z,�x�j�:M�C�ʛ�mf�5
���cu��ޏ��!Ɯ�J�9e{��b*�*.| w���6�T�=�|��M�|�$���(�����~�^�7~�z{�#� p%��t$]-!�r��|&�}��a���Oh%��|w'�ٟLgi�R�,�4[v�LGI���N���O�=]�7����@���k���X������I�KK�hD�6}_���	��@5������1FP�N3O/84��1:ߛ�?�KF��� {x_S�x�����1k��&ط�+D?���~�3��P��Sg���F1�@�:��1�Խ ��j��5����qG+�TS��Ȱ�@�{�h�e�д�Q���@wam������G���hV�w]�;��é��HlSX���c8���k\�\Թ�X��� ��"\�ݿ���\jF�d��D��rb���E�:�ǖ$�RŤw�]Z#UıI��HbFcg
�ö}y���\�*�[4��N3H�;G��)[����h�w���DsG���Gs���9�':����ꢶ�t��n�v��e�9�J�_���@Jt���1&E��vE���!d|Fg9��Q���Ě��r��;��^@���� x6�s��W�9t�ԷpB�{��j��t��m�ϧSc�PA��C��!�v���fC��&�%��o�D g��e�rYۺ4o�-�7q��^�G�^k�4>��v���T	�|`�$�1�=�-oJ?�I��S4��tգ��U��<H,�� @ �oG��d0���~�(���+������������"Y���{��z�]0l*v/�6~�F����ix�������J��^�[l ��CC,���S�;���r�,�X>߹������;�	\f�ṑ
�R�u��=p���(�<���c}`�*ag��5cT�u;�M�9Rd�/���k���s*�@	1��S{U6��}Xr��S�nSġ�h[�]��txrd�U�ײ�"1�G�^����.�"�0���6�"�JMy���:m;�q��-<|h�̖Bd�oЕ�;��Xz�?���{N7ڡ��ly��5��å�$�/��ޓ�]9&�]H��\��evn���y."ˏ��DO:lߒ�׳���R�,��^0�}��o���9�7E@��O,i���xtesK��xE�=��)���ʱ@[�`�OL@��'�FR0�ja����`����@�M�o�s��n��������
��6n�MF;.]	N�;�@@��p�{�P'd��G�e�#1��t�W&{�Zx\��?=E��;�0}_�! �WL�^obB>�z� Pr)�d�F-�>M��hs.�\�ڳz�wO��ԯ�����h#�I��0�F���M>�s�h���h �\�C1�yd����p�L��j��9�w+Ro�`��hZ�T#2}��ޔG!��5�]�,|�Pvt�yu�b�DH5�2��3������$�`�#x��E\ؑ�r��y�x�k����Fq��(���+�˗I�YM`�f
��<�f�= ���|H�����(T<2���H"Dt����wP����W"U߬��������w��	D�E5�|��S�H˪�ђ緾��!^h�%��35P8�؜�9ɾ�\��~�䅘�0���t�{��_%4�=���-8�&>�-Y{�V <'�'��u���dMu
�a0��=��Z�`਍c�N2veq���"��Q�;��c�S�6��1��z��2�����΂-�;�ȴ�fr�W�ʳ�GG���ENkUu���晑��)�dj�F�X�)�@y�`f��2S�=���pJ��M�)R�մ�Ǯ�6�
����=�iw���`�d���q�I�lC�Ss�9�J�Q��px�t5��,�����#x9o��J�Ʀ�e@�iOK|!~�5���aêj:�\O��6Ć:�I=#0A�wO�Z���P����ћD{$Ti�'_�̶eB��^?-�Ӧm#�n��oRª�(�kt��X�b�|J�:���8V�3��1�d�@E�=�5�m��4*2;�^�(]��x��X��������G�8A�B7�.�k�᧴5lb,Ɣl�%qӤn���\��_0P���}��5�``!w'W`��H�0cae�<��@������a�cR�T|�<4�홌+��ݴ��1��*ײG��-���ɇۈ4���L#�}�������R(������j>q�t�*��J�"��������-3�K��VO�`�)F��PߌT��^*������"�+�Z��nh�ڱ�Xk=*���hb6�L���Q��SVt,P�9�B=�2�v_�\\o0�(󂂍ղ��@��U^-?��&_�p�a��9��M����cRv����o5R:�|u�`�`doͶ��6K���@n��$��;g����ܞ���6F���|�qx{;k�Xm��)Z�SXʢ�AR�'c��)( 候�J���غr%	�W������y��ȣ��yG�iH�ޏ��c{}����/>��W߯�K��*T��qt_���n.=�£o�x�c~�� s-_��<�%d��Yi�չ3��Z����7ᆞ|��L��������&tC_C�uA�ߎ%��F��}k�zZ�����A�*��x�K?�Jw˥�'��g��'��j��������P��|�Fҁ9ҺdN�y�P}�<_h��4,��d�����_��ދ������!A�)�_�oD�xso�6ว91�����[�*�6����V��<[S&{��&�Ibg;�׺��&$?�_t�����ѫ�|���*ʤ�.�bɸ�$�vʴf~�\Ǐ��9z��D/�k,�����	�8g7�4 �<�}��>�47w�K��ے��P�D���}ǐ��t`�����mQ�FG��V���y)y��'��ζ�a�ߏ�R���a�2��'���Z6����Τ�)�}�x�<�%�ߏ��6�{�mЩ�ت�<��cŽ|"_<��W�����Q��`�C���L�������Wdج���8�A�u�MY������yr�K�e ���i]�)��Y�I�F��W�'#�|��%N�- ��hb+��#��w�����\K�\W�b%��{�)�[������*h�R�m*W&���٬�+/h�r��P��qr�{�j�A��zޫj���[�����	 ���}%H~81����tdw_D#Ů��\I�\��O $�0�EF�k_�P����j��D<|�ں�t��Rr�β��W)��.B���&�NcC���Ҥ�s�M�k�����,!9:ٔBjaj�
�E2lw�D"F1��r�6�Rt�tf�\����Fi��}uV��$�S�ob�6��yL����-�!�?z�o{JL.��ӻ���N��	E�E���SS����W�2p�vb*��y��-O��Cv�&Be�ѫ�Kz�)N]�m�>,m��61�_�;��2�ǂ#:q.�Y]��\+҄�~��ldP�0m���e{��gҦ�N�:�>�MՇ_Q��²�,BC,���A�������+,���s�&��ZN����ⅉ벃�d���T�8ʐ��5�i*��cT_��#tވ�=T��Qt	��]�}��؉f��kǑ�Te������Y���6�5�V�Mj{��*���?���%x�J5Ǝ� ��"�{?ԫ>���(�t�2ϟ�5!cL��?�+J�J���ȝ^���<�Yc�����+�O���$�|z�ڣ�IMFv�a���7�;�J[���;�N�#>��w��|�g����e	�`^���l,�3a"�ڧ_@��J�&E�H�1��i(Z�g����ܝG3���-]Я�p�h���ѥZdMz��o�K��]����h��'P�ܗ��T��.(�˺T�:z�CU��慴�Cұz�4�f1�ցk
�G1� Ӻe"M� �¯;ٖ�\��ÃM�8Kj�'�k�G7r4D!��=�K��9#�^���'	�=b��7O_��\��?J�S�B��/p8�yZ�1��uG�k�J@�i�s��륶��N�3+�`v�A/S^�+�,N��[��|'���P�����l��Pφ]�l�~���DH�M��׋�����D�>���&�LsWhs{Z�Q��P�L�,c��*�t�M~Z�ћ�"����9�~����� 1,�����0:>^^� 6z��O�{�Rq���2�e�6����jC�`�E��wN|�}����°Ft8~��Nj��؍���4�q��5	�	��$HK[bR�e�-����iwOw=��SAa�	�`������:j� co�]�჎��WV�O�	�C����Q�Ky�KC��p�L��-�'�o]u�9)b���Ȩ�ȁĿ1{9?�`�,���@S)��u]�T�a[��Ņa�|����!��5�r���n���H�,�#�t^��u�'���� 0a��`͉*�"'뮡{L��*�ʺ�>1�&��Kk����<.�8���9���<L{�P?��x7��D��|�l�Rxh~�����[!ۑk��[����4��l$��;J�^"�D7�	�y5���^�&#ٖH�u��16��+#�&t�/)QV��b��>�6PH��nr��KI	�-R�|t�I+**c������۰a=AH*�؍�<yA��E4��-�u������,R
!��V��'�V�u�9����۽ŵ�8�-{qgJ�Д��䫽��N���?|?*�i�|*�s��	�: :�w^��9W �\���aL|��ߌ[��3��L�1¯�ʬQU�K�ԥ4�����a��TX���|��@�8��έe�⋿Ax�:�;��vc�%0/�D1�I���f��
���[�m�i"tR�)��|��.���arr�"=�`�� o�W?}��Ø��	]c�.��5�ZH�r�A������9�8��D�Kؓ���ϘV?���<����X��pG-��W��{*j�V�Q`��{�J{�P�/��zE��^���m�Y���V���Y%/��û����"<�[�%�_	ؖQo�옯�T��i� x����ʙ(ǩ��a���]��6>s�ţ!|�ʊ�x��yn$H�F��! p�[���G�k�x+
M�S[�@���
ѽT��T��}�!�J�Bivm�·��0~���D�`���=.�R� ���|:�)��Eƛ߷2�<�9�3@��A��΢�^ ����<��ETZ܂� �w[!:�)6W�$?���#��\_sĪ�t?0���&��	�Y�ޟ�H�vQ}'b����x�qD�KJ���8�f��L�j����ylgNb�"��k��d�f�)x��ʦ��q����	uÖ��]8�:͟*)5�#�{vO#�[�϶Z�vc�U54�!붯�M�]b��d+��,@�S��������HH?�i�?�q_�IO\I�g��Uj��V�Hf�o��<� �Ҽ@ɂtPr��X)P;��>�?0<.4���v�G��_���>WCã�W�w��s�BaM�²w�	�n���L�7<�.�)u�zAP���������Ft��ƞz�6���O8�:C�-�uA��������ܖ�G�6�q�&*�lXG�R�^�Ap�@j�f��C��F^=`�尙�9B놳���]D����U�sC�h��Ƚ��d��[�����琇��:��ۅ'"�9M�&ߩ�9���T���s稴]0ވ����gV��!�4�������g����Su�	����V��vv��7��=E���7��q����0����%B��E$Ip�||��(y�F����{ �[X8�ws+��t{�����l��L�=X��	�Ln.$��m	��xEl�]���?��3�X��l��� ���T��oӞ��㏳(��7Ӟ��;(f��wg#� ���a�Q�ק�~i�~� ��!��P6�U���B�M�m���c��0R����:	�����}�tH��$*���}p�c'����O�a�a��� ��p��j>$� ���.����^�8�7����F%G�9A�)]�BB>���|Ϳ�?5X
eb�pI1���\��F֭+ ���8򃏯�2�#����t�U�����������#��舖ժ��ON:�eFgs