XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������������[/�C���n˜z�,�MZf��q��ަ��h|�iǑ �{��\�����oɌ�e���K��ʶj�ظ�8�G�7�\m�a�G�j�v��;�U&x�d:��}��dy���ٳ�y}��7����9�n���a���ro�����Cp���.P��KHc�ӭoa@�N�z��C�ˀP���=�u�V_1�����9ķ��@�~&@�D�iZb
���X���j��"�F#țK�N�^�׀�0�rc�_U`eK"p=��]>���Λ�iȧ@@Ve�n�2����Q=�Kі^T�VO���B^�����aC*�֋D�;/kS�?��y�f�:�m�de(Lt�!
��h%�V��� %B����쳺��}�R~EἀV�L�W3.�z��5�	i��Hv^�ӻ��A1�X���K�<�~���<,a���_��)t:��c�Y>;1��g){}8�V׳���%�k�6�z�x?�uxeO��U�J�˟[ܶg��&ǩ'J��zf!��vd۔Ѳ��䪩������_Ą9]��`C�����+c�d/��,�#��K��gVɻ��A�&_�l���y^$�όd�,�M����W)
��{F�}{�g��6!�N��Ǌ}����Qv�
s� �b!Co���}�b3c��K��~��x�)ɗ��/ ج��t�mc i��vE{�%���X��{��|�棇�BR����c��Tz�pH�����~mq���ow�J��X�oć96C��;XlxVHYEB    dd8f    2160V�Y�%�J��1�X��i��� Js�F�����N�J��ƜfK/	~A����\=Y$%�L�I6�h�\�"!aQ(�C��i��9�N�Y�L�S���M �h�`x�V)ڿ�K�����u�C����}o╥hd���� �wVNj<�����_Xa'|>(��0�|�Z�8�;��1����(���R���W�B=�P�+��&��-+K�@�"��2|���m�17s�� Z�8��:��=*M�H(��5kS�X����Ȭ�b�je�ۆE��kҸ�U��,o����-	4P�i�l�I�;L�_f�2	S�Y�;3&_P@�@9����x@��A�،��=��M��&Lc\<��W3���{��AV��;�Zh�U�3�u�X?�^in����Ҽ�5�h0�Lx%[���,̋���2���v��i-���V�8�e�������Ҷ0Uf���4:v.��ڵ�ȵ���[������L�O��Ơ��qUt�c,yU��+��@j'���?��Ɛ}�A�ZX2#���A����� ��v8M�ZfR(bJQS�P^d�9�l���+C"�~(8_�"-}�E��&&�=�"(`0	�m�I���n��O翦z�LCK���~ך��Ll��W^?���/��gk��!N]øe��!�oiXQ��1�����;�=���3��)���z��~���
��=���hWX�w����#��f���)o��ܝںb�ݧʅ��ڗpD$�x�}
;���A{���횫��o�=��Mz'>��Z�Z]��UX'�3-'_1d�������οN��&؇�t3xp
�+.�LC�\�y�t��J�+L�z��])�D�QN,��u���Z�wߗxx@��;w����1Vmq�WZ)��a��,V�֢�d~��Ҽ!8>�\X6����j��%��-OΕ�RXu:(����9~
�LBۂO���c��i��V(Z�͔/޶�6��K�a/^�4����o����Sy�0U����NZ~��?�#�k=漚j ,�R!̞��<��
rv��?� 4����b�cQ����}��9��@$4d.L�j�_�(ϓ1�BU���"	=�V%��5�N�8�y�J`ۨǡ=q|r��+0l�K%Q�.� L�2B-�
�|YL�x�Qz�q�9JrI�:�/{������W�ɞG�ފI����V��P޴��)V�������$.���4b��q�'�,����T��D�����#�:�	X�y5d-PwQ0hH��p�(�a��t�N��v��9��	��X#�A���ahg�ꁓ��ۙ~�vr��c�9Z$�t�o�{��0�����.�'N�tcD��Rn�k̟K��Yg�B~�%׏*�_|[�~�jiL&~�Rf�y�>!֓t���N��M}?�tG/��o�KT�$!-"Z�I���Y���|���z�c*���fR�˫4�̯ ��t�~z�T/��`U�-Ix�m�%��p�v�\���⌮c�����01�a�o�f�`@Od��cꑖEǳ���Y�W��AKi�`ѲET�T4>��T�K�/#�?��� \,�Zt�駺��7���E��9�h�h�e�gs�\4�h���
^:&-�ϢL :���s����~�A�X5\��ۜ��:���.0k�r��!�=�1�	��ř����$ݠ�L)i(������*�^|-u%$��Dp6V::�IF%tt�Ҕc}�(��Dn��o��[ȨJ&�e{�,��)m��t�������`�n:�i��"���8l��Rc w?�;��9�'��dq<�6�4���	�vᎽ<�G���p��M�c����6k5%���*e�)B��r!`��uM���#��'f��`\b1�71������	C�F�?K��y�����Z��)(FN$��N���L�>�圫�p-��:�Ѣy*��l�$ο4�O���U��i��	�p��:y�#Z��P*��e�-҇$�����Z7%� ��*�u�H�K�6�?W2��T����D�q ����~�*N�U
]��s}�f������o�k� ��n�mKܕ��� e����������/B:jL�'А�&�53��qU�I۾�I��PޒX$#?n5�/j�[�rjeS��<�fE�`���@�/?�~8�N:U��<d=q��|�:[d��V��ߧ�L�M1�c��j�DE?8�e*��G�ӐM=��\��'9��gΌ���v�H����wV�8N��ck>&�Y��2nþf8��b!��e�Q�_x+`�v`A�����Q��)B`�d��(=K"?c�8�@�����#�ї��~�9 ���>���O����.V�㲹sT[���n��9��~;��#���y��P�����L3�;�n_ ��"R>j����v��xC���$f+y��H"\Ҵ7�C�!�Oh��(�.>4�U�!)�=�ٴq���N�Ԑ:gS�%��E�d��Im������ t�Am&�VR��Jy��b�ߤz^��Ek�O�h2�?�����H�C� V~b ˝	���}'3I��,�#2�{Dl ���bM�h��p�����72��iJ��<�%Z���Ⱞ ���ˆ�����~Cm�^'X0x������"�Z���X�D����0�	!3�T���'��o(�h��a��+��+ܽ&�`���&S�� �ϡh�'|$_�ϐ�6͜J��)D��o��������ە��tD�#���SR��)�ce��
�g�S�_�'���2v�������>���+*@���r๔i��5�iG���Q�N�����T�
N��@��s��c�xCV3"����n��/�(�[h���󬍓H��q��hk�>�=!L��_�tD�y������0Ji*}��އ�KN.��LjZ"���G
��|�3����:�N�t�҄����sM�[�t\/���:h�ϊ�L�3�<DC}D��p[Q�T��K��BX����fw�*y[��ɒ>OF:o��	����^TOJ>�]K+���hjЋ��'�R��hd�������ʌ���zr�c,'Dbʠߑ֦�'@V�rc�NϚ/���݀��h��2�ח��	�G*Q%���M���?��)	�?��5�}oc�hH�8�Q��L������E�k�%f`�t{h���o�+�ϙ��Jt.��ݾ+5r�p��N���H_�iUs|�N���L ��˂�py2G��a�n�_HƋ�E������a����̈́��y�X3v���x���x��(I�]By���A/��#�M6�{�:���)��Vm�,"���\�8$��a � ���u���Z��fj#���Q1:��3�u��|���/�"�bS"�<�h��	�B H�4~�f �'P@���������GW��	�Z	B��g	
�2I�\T�(�޽���6�OҸ�����/t��	{%��l��f;3�g�
�`�ݷ���M7ゼY������I��8��:��b�K���֙v(y���r�ٯ���o�"��e9����zk���PDv���D{�Xŵ�qIt� ;��)A��>U��e�`�1]� w��)�F,��:����o�sfk�-L�\�n��_mj`C	�IH#J�����ۇ��al'09(ΐ��x4�T5ʆb�Qꦍ�WyF��YQ�S�q�?�5¡x�k��5��'dV�H�@Yd#%q�:����$�_D����~ƴ���
2զ�29���R�)o;��ALi[���`�����F����}�%*L��� ��]��0g�ឦU�UÈ�8��sE���U.Y�����|h���>'���%O��p������'�) ˴c�M�bό�����Whp5��<�gM��O{>���;�� ��g�9a�^�`ʪ��U!�6 i�]`,=;.v�ᆊ�H�q� �~+Qh:L%�Ϣ>]�3gV�ˮE�Z�� ���Č�#!�D����#�o1;c�ZbO�Ve��(T�>q��fY���i�/8�<��E���oi�z�D˭^C;��zC�&O�2��$�Dv�)@��Łw��x��Fȭ�'�Q}�r�L��e� �<f|Ţ#�;�۫�8+��,��񑹸y�)��v!&����4zO
B�~���j��f�fj�n2N-ǈ�a�p5�=l/_ ��Ԥ��M�T�����Ǥc�6N���C���Bvhȧ�0�=^��^��I��sn�G�x�o�My�W]���a����J���*�S�$�_����auךVp-Ģ�I�c���'vN��T��ȋ��:e�5��u�*��X^wkR�-�St��h7�ZAJ��M]��9aW�c�Ϯ�9���y�cʘ����5b����F剱�C�(Є��p�Q+����ͳ�E��ڇiEPWA:��D��G"P�N�ɾ�vd�c��u�9d�c�w��b�,qN�'9�����T�RR��N-{��'aլ�9X>��eR ���i�'��0����+�`�*��B�Ўʬ��w?�Һ�w�%S�(��jRVj�D���]& ֤�苜��ه���)T���2�+�9���d�j��9�s{��ظY�\��s �����%�!�&n9�bz���]砵*n���-G����U5�E3u�jMnw܁LW-��(N%/�.fm������v��;�
�G=�y5+kb�蛾�ڒ��U��� ���}+p���a���:Wf�&���2�}Z]������+~"+%M"�%�/?W|�5=3�QBP�m�Lp�dܻo�����I&��7���$��ZH�;_6�HC<I�B~!��>�/��;�,�,T�����
m|��9(3�A1>�Sͺ<b�4�:_�C��>i��зA����u��ab��J�"(	��W�gnw�����А�0Yl�i�.�B�L�J��2��sa�gҘKh,������?b+��ˈ{ �5 �݀|)h�Q��*+��4U �^~6 !�lp�^+�m裧.��L������5k9;�#�F�{:�0�`q�%7���k��	�d�����a�4Znq�u�t��Mbx6��]�g�;ʣMm���;dO��5i�
��v�NJ=���<�(��P:��ŵ�G_���~HUk0C�fKS��
/C%�-d���@��R��t�TG�������T5��A]���o�S�.'�6���X	j�)���*J.�S�a1�� �=Q#ӌB	���K���U105"2Vds@�P���U�G�OvJ��E��;�p�I�З�8�΅�������V�[�1�9�.�}^xT$�E�O+d~j�KQ�k���=��fz�駊_�|6�|��`К*?��|��Vw[�e�xT��M:8��`pM�y�5���LO&�u�J���0�w�\��W[qݪ:�u��Ĺ,0y@{d�R�Mp4'0��W	'�W����X�Y4� ��cm̖����ҷ��\���3 ��?�³r^���ӑ����_�>�O���J�鷭��+>�_����Ž��q�i6r�>B���ߘF.�TL��=�F\��aMT��l��Cz��A�ֱ�̫���+4��.S�N~��2�[���۰� !���`n.FSy9�sk�x1����՘�:�r��O\#�	%4@}�y|�]���1�-��X�r���݄A1��JQ/�i����Ŵ�	�����v� K!�T0��ʺ�2I.2-\b�b�q�\��w[�e��g˔{�|q�tX��)�B��7۲�����-f�QI�i�p�v�L�6�h���=F���x�糿o���U��7pS�v�W%�ұ�r���?�'O�٪0߫V�Mp^+k���ӌ��,rs*_�+��d�.�4��l���Ly�[�!�/��<f�Ii�Z5�&��hk���a�(�rG\�H�w����]G�V�<�FK̝yD�6;��������߸�7����o0��
��b��W<O
5͢�RL��V	�}�hZ��ZK<���߅��|���L��۟��SQ�U\Ŝ<��-��J�6�/fv��T�5��L
g����^}�� 4�a��]×-@�����7Sz�qr��><�m�b�m�r3�E�!%�݇:�C�:{����;�.|��WL�:7u�f�C}t��o'qZn]K�	�fF����"qՎ�ڭ8.j����[�M�C��h5�3K1P�N �N��Tϵ%��I�y��Y�wI��JV[Qg���ђ*�P��s?�����&L��6�q��j��}�f�7�����;6����:#�8�O8[�S�PM,�P%�j�t}_A2�-�Xa4��o���ڛ\S=���ɛ�]��K�>��%��j�^�~���b��$��d5CV�J���q]9����X���9���Q�2�N"D�[d��8�(�(z�p�Z(]�v�3���H�fc�vr�	���C��t`��|��H��-N�N��%ae�_9����ȊD��uX�x��5�sI���d�C%< �56�`�4Q�a���� L(p�}Z»�7Z����H��0�r�e��3�%4<��_]:}�#��AH��m��U�]��Ly��לΚ՛�i�
�oH~%���i���lp��!��H/`��H��ޖU��o.���
u�ҋn,ycmL��5Ϻ�r������	�@� �j��A|�� �{���d����:�,)v-�=У�ܒq+��31�CN��Y9kc��?�&����Iz�.{����`0��2*�B.���Ӌ��*� OB���X�����'zT��U�v�������h�60�����K�A�F;�(6�(�}HV�N��c���}��,��ڎR}��&�ٺh$�ti�ԋ�9��	^Ƽ�b�% ���Գ��#�h��zC ���P��JY͘�O��d}v�S9m������Ø��yaaj+0m�b�7yT3�B�҅̈́ҪB��!u�cbG�,�T���b�����;u��Is��BJ���������t�Z�"W�WH4_}�����v���KhR[�u����E�
�>(OVnd/�;�S ����oM�*��!B#yH?�E��1�OuHTqs�T0P�O4����c���%F|l5Ao�<k�*��T�Qw��.����"�!�9�5RDz/���#p��Z_�l_��*s�,�Zo;�ż����d��O���yMH�"�$J
���\���̺>�E���n\���5T��L�n�I��Z6���爔�i�g)��h���4�l����*@�ނ��v�������?���'�12�v��$�At]��7Ƌ>N����b®�&㟙�����-	�d��@�0�)AEl��I��64��;h$F%	�O���91c�wQ��ҽ��\t�CR��0͇�2&����Mec����Bg���9��8� �+q���@�c���䛡�����{�� z!o#z�c���Fɬ�G����?��?	P�����;8�+��S^Meg����W'���ۢ�@�	��ٓ�ma-�&h��Pm�,��L�Z(�X�Y=�L�cY�����NWys9b�������2h·#��O�lG��	uDF �����V��[�����>v) ���R�Ŋ���Ѷ:X~��>^�]��Ӥ0�����r
��_��N�l`+C���'w�9%(�'Q�,n�kV*��:=0^�����Q>��oZ���>����!�V���Q������㩆{�Қy�L���-f1��U]/VB�M�]��}ng1��ǖ�� �� �'1^|5�Io��@m�y�E����1Qu7�۔�|���a�y��$���2aЊ6}�� �v7{b��!0 �����c>'t�e�3��2���%A�b1 3~�����J��_�p�X~�O����^|Sd��d�n�2�.��!4�K����Ɠ�H����Y��9q�\�j@{Q�M��r4��őX�����K��6IZ�7$��3��ux�?�,�4�c���K�r��\�w((����b����ګO��K3�f{���+�/��r�K�&"]����R �e���AUH�n�9�P�y"/S?W�]���/�������@K���s��f�������h���4��g���HjK��8�_���,��`$�E"�Y���"��z&C���Ů�b�_)цW���A��?�l��!�U��u� �n�}�M®����]��Gp�'��fP/E$k��5r�C�ב��˩��m�T�`8��Y_����������Y䗅g�|�<+�(U�AW֞5��ުv���+�ަ��0�������� ��ܳhi^��p�;ǲ|#��Ï\(~�8M�3�>忘%]�[�QQh4=$#|[�ҝ�����A/��4�a�E�}&���n?u0�))��^��Z�	࡙}���Q�#K����i