//-----------------------------------------------------------------------------
// system_processing_system7_0_wrapper.v
//-----------------------------------------------------------------------------

(* x_core_info = "processing_system7_v4_03_a" *)
(* CORE_GENERATION_INFO = "processing_system7_0,processing_system7,{C_ENET0_PERIPHERAL_ENABLE = 1,C_USB0_PERIPHERAL_ENABLE = 1,C_QSPI_PERIPHERAL_ENABLE = 1,C_DDR_V4.00.A_C_S_AXI_HP3_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP2_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP1_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP0_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP3_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP2_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP1_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP0_HIGHADDR = 0x3FFFFFFF,C_GPIO_PERIPHERAL_ENABLE = 1,C_GPIO_V2.00.A_C_EN_EMIO_GPIO = 0,C:GPIO_EMIO_GPIO_WIDTH = 64,C_CAN_PERIPHERAL_FREQMHZ = 100,C_FPGA3_PERIPHERAL_FREQMHZ = 25.000000,C_FPGA0_PERIPHERAL_FREQMHZ = 100.000000,C_PRESET_GLOBAL_DEFAULT = powerup,C_FPGA1_PERIPHERAL_FREQMHZ = 150.000000,C_PRESET_GLOBAL_CONFIG = Default,C_PRESET_FPGA_SPEED = -1,C_PRESET_FPGA_PARTNUMBER = xc7z020clg484-1,C_SD0_PERIPHERAL_ENABLE = 1,C_UART1_PERIPHERAL_ENABLE = 1}" *)
module system_processing_system7_0_wrapper
  (
    CAN0_PHY_TX,
    CAN0_PHY_RX,
    CAN1_PHY_TX,
    CAN1_PHY_RX,
    ENET0_GMII_TX_EN,
    ENET0_GMII_TX_ER,
    ENET0_MDIO_MDC,
    ENET0_MDIO_O,
    ENET0_MDIO_T,
    ENET0_PTP_DELAY_REQ_RX,
    ENET0_PTP_DELAY_REQ_TX,
    ENET0_PTP_PDELAY_REQ_RX,
    ENET0_PTP_PDELAY_REQ_TX,
    ENET0_PTP_PDELAY_RESP_RX,
    ENET0_PTP_PDELAY_RESP_TX,
    ENET0_PTP_SYNC_FRAME_RX,
    ENET0_PTP_SYNC_FRAME_TX,
    ENET0_SOF_RX,
    ENET0_SOF_TX,
    ENET0_GMII_TXD,
    ENET0_GMII_COL,
    ENET0_GMII_CRS,
    ENET0_EXT_INTIN,
    ENET0_GMII_RX_CLK,
    ENET0_GMII_RX_DV,
    ENET0_GMII_RX_ER,
    ENET0_GMII_TX_CLK,
    ENET0_MDIO_I,
    ENET0_GMII_RXD,
    ENET1_GMII_TX_EN,
    ENET1_GMII_TX_ER,
    ENET1_MDIO_MDC,
    ENET1_MDIO_O,
    ENET1_MDIO_T,
    ENET1_PTP_DELAY_REQ_RX,
    ENET1_PTP_DELAY_REQ_TX,
    ENET1_PTP_PDELAY_REQ_RX,
    ENET1_PTP_PDELAY_REQ_TX,
    ENET1_PTP_PDELAY_RESP_RX,
    ENET1_PTP_PDELAY_RESP_TX,
    ENET1_PTP_SYNC_FRAME_RX,
    ENET1_PTP_SYNC_FRAME_TX,
    ENET1_SOF_RX,
    ENET1_SOF_TX,
    ENET1_GMII_TXD,
    ENET1_GMII_COL,
    ENET1_GMII_CRS,
    ENET1_EXT_INTIN,
    ENET1_GMII_RX_CLK,
    ENET1_GMII_RX_DV,
    ENET1_GMII_RX_ER,
    ENET1_GMII_TX_CLK,
    ENET1_MDIO_I,
    ENET1_GMII_RXD,
    GPIO_I,
    GPIO_O,
    GPIO_T,
    I2C0_SDA_I,
    I2C0_SDA_O,
    I2C0_SDA_T,
    I2C0_SCL_I,
    I2C0_SCL_O,
    I2C0_SCL_T,
    I2C1_SDA_I,
    I2C1_SDA_O,
    I2C1_SDA_T,
    I2C1_SCL_I,
    I2C1_SCL_O,
    I2C1_SCL_T,
    PJTAG_TCK,
    PJTAG_TMS,
    PJTAG_TD_I,
    PJTAG_TD_T,
    PJTAG_TD_O,
    SDIO0_CLK,
    SDIO0_CLK_FB,
    SDIO0_CMD_O,
    SDIO0_CMD_I,
    SDIO0_CMD_T,
    SDIO0_DATA_I,
    SDIO0_DATA_O,
    SDIO0_DATA_T,
    SDIO0_LED,
    SDIO0_CDN,
    SDIO0_WP,
    SDIO0_BUSPOW,
    SDIO0_BUSVOLT,
    SDIO1_CLK,
    SDIO1_CLK_FB,
    SDIO1_CMD_O,
    SDIO1_CMD_I,
    SDIO1_CMD_T,
    SDIO1_DATA_I,
    SDIO1_DATA_O,
    SDIO1_DATA_T,
    SDIO1_LED,
    SDIO1_CDN,
    SDIO1_WP,
    SDIO1_BUSPOW,
    SDIO1_BUSVOLT,
    SPI0_SCLK_I,
    SPI0_SCLK_O,
    SPI0_SCLK_T,
    SPI0_MOSI_I,
    SPI0_MOSI_O,
    SPI0_MOSI_T,
    SPI0_MISO_I,
    SPI0_MISO_O,
    SPI0_MISO_T,
    SPI0_SS_I,
    SPI0_SS_O,
    SPI0_SS1_O,
    SPI0_SS2_O,
    SPI0_SS_T,
    SPI1_SCLK_I,
    SPI1_SCLK_O,
    SPI1_SCLK_T,
    SPI1_MOSI_I,
    SPI1_MOSI_O,
    SPI1_MOSI_T,
    SPI1_MISO_I,
    SPI1_MISO_O,
    SPI1_MISO_T,
    SPI1_SS_I,
    SPI1_SS_O,
    SPI1_SS1_O,
    SPI1_SS2_O,
    SPI1_SS_T,
    UART0_DTRN,
    UART0_RTSN,
    UART0_TX,
    UART0_CTSN,
    UART0_DCDN,
    UART0_DSRN,
    UART0_RIN,
    UART0_RX,
    UART1_DTRN,
    UART1_RTSN,
    UART1_TX,
    UART1_CTSN,
    UART1_DCDN,
    UART1_DSRN,
    UART1_RIN,
    UART1_RX,
    TTC0_WAVE0_OUT,
    TTC0_WAVE1_OUT,
    TTC0_WAVE2_OUT,
    TTC0_CLK0_IN,
    TTC0_CLK1_IN,
    TTC0_CLK2_IN,
    TTC1_WAVE0_OUT,
    TTC1_WAVE1_OUT,
    TTC1_WAVE2_OUT,
    TTC1_CLK0_IN,
    TTC1_CLK1_IN,
    TTC1_CLK2_IN,
    WDT_CLK_IN,
    WDT_RST_OUT,
    TRACE_CLK,
    TRACE_CTL,
    TRACE_DATA,
    USB0_PORT_INDCTL,
    USB1_PORT_INDCTL,
    USB0_VBUS_PWRSELECT,
    USB1_VBUS_PWRSELECT,
    USB0_VBUS_PWRFAULT,
    USB1_VBUS_PWRFAULT,
    SRAM_INTIN,
    M_AXI_GP0_ARESETN,
    M_AXI_GP0_ARVALID,
    M_AXI_GP0_AWVALID,
    M_AXI_GP0_BREADY,
    M_AXI_GP0_RREADY,
    M_AXI_GP0_WLAST,
    M_AXI_GP0_WVALID,
    M_AXI_GP0_ARID,
    M_AXI_GP0_AWID,
    M_AXI_GP0_WID,
    M_AXI_GP0_ARBURST,
    M_AXI_GP0_ARLOCK,
    M_AXI_GP0_ARSIZE,
    M_AXI_GP0_AWBURST,
    M_AXI_GP0_AWLOCK,
    M_AXI_GP0_AWSIZE,
    M_AXI_GP0_ARPROT,
    M_AXI_GP0_AWPROT,
    M_AXI_GP0_ARADDR,
    M_AXI_GP0_AWADDR,
    M_AXI_GP0_WDATA,
    M_AXI_GP0_ARCACHE,
    M_AXI_GP0_ARLEN,
    M_AXI_GP0_ARQOS,
    M_AXI_GP0_AWCACHE,
    M_AXI_GP0_AWLEN,
    M_AXI_GP0_AWQOS,
    M_AXI_GP0_WSTRB,
    M_AXI_GP0_ACLK,
    M_AXI_GP0_ARREADY,
    M_AXI_GP0_AWREADY,
    M_AXI_GP0_BVALID,
    M_AXI_GP0_RLAST,
    M_AXI_GP0_RVALID,
    M_AXI_GP0_WREADY,
    M_AXI_GP0_BID,
    M_AXI_GP0_RID,
    M_AXI_GP0_BRESP,
    M_AXI_GP0_RRESP,
    M_AXI_GP0_RDATA,
    M_AXI_GP1_ARESETN,
    M_AXI_GP1_ARVALID,
    M_AXI_GP1_AWVALID,
    M_AXI_GP1_BREADY,
    M_AXI_GP1_RREADY,
    M_AXI_GP1_WLAST,
    M_AXI_GP1_WVALID,
    M_AXI_GP1_ARID,
    M_AXI_GP1_AWID,
    M_AXI_GP1_WID,
    M_AXI_GP1_ARBURST,
    M_AXI_GP1_ARLOCK,
    M_AXI_GP1_ARSIZE,
    M_AXI_GP1_AWBURST,
    M_AXI_GP1_AWLOCK,
    M_AXI_GP1_AWSIZE,
    M_AXI_GP1_ARPROT,
    M_AXI_GP1_AWPROT,
    M_AXI_GP1_ARADDR,
    M_AXI_GP1_AWADDR,
    M_AXI_GP1_WDATA,
    M_AXI_GP1_ARCACHE,
    M_AXI_GP1_ARLEN,
    M_AXI_GP1_ARQOS,
    M_AXI_GP1_AWCACHE,
    M_AXI_GP1_AWLEN,
    M_AXI_GP1_AWQOS,
    M_AXI_GP1_WSTRB,
    M_AXI_GP1_ACLK,
    M_AXI_GP1_ARREADY,
    M_AXI_GP1_AWREADY,
    M_AXI_GP1_BVALID,
    M_AXI_GP1_RLAST,
    M_AXI_GP1_RVALID,
    M_AXI_GP1_WREADY,
    M_AXI_GP1_BID,
    M_AXI_GP1_RID,
    M_AXI_GP1_BRESP,
    M_AXI_GP1_RRESP,
    M_AXI_GP1_RDATA,
    S_AXI_GP0_ARESETN,
    S_AXI_GP0_ARREADY,
    S_AXI_GP0_AWREADY,
    S_AXI_GP0_BVALID,
    S_AXI_GP0_RLAST,
    S_AXI_GP0_RVALID,
    S_AXI_GP0_WREADY,
    S_AXI_GP0_BRESP,
    S_AXI_GP0_RRESP,
    S_AXI_GP0_RDATA,
    S_AXI_GP0_BID,
    S_AXI_GP0_RID,
    S_AXI_GP0_ACLK,
    S_AXI_GP0_ARVALID,
    S_AXI_GP0_AWVALID,
    S_AXI_GP0_BREADY,
    S_AXI_GP0_RREADY,
    S_AXI_GP0_WLAST,
    S_AXI_GP0_WVALID,
    S_AXI_GP0_ARBURST,
    S_AXI_GP0_ARLOCK,
    S_AXI_GP0_ARSIZE,
    S_AXI_GP0_AWBURST,
    S_AXI_GP0_AWLOCK,
    S_AXI_GP0_AWSIZE,
    S_AXI_GP0_ARPROT,
    S_AXI_GP0_AWPROT,
    S_AXI_GP0_ARADDR,
    S_AXI_GP0_AWADDR,
    S_AXI_GP0_WDATA,
    S_AXI_GP0_ARCACHE,
    S_AXI_GP0_ARLEN,
    S_AXI_GP0_ARQOS,
    S_AXI_GP0_AWCACHE,
    S_AXI_GP0_AWLEN,
    S_AXI_GP0_AWQOS,
    S_AXI_GP0_WSTRB,
    S_AXI_GP0_ARID,
    S_AXI_GP0_AWID,
    S_AXI_GP0_WID,
    S_AXI_GP1_ARESETN,
    S_AXI_GP1_ARREADY,
    S_AXI_GP1_AWREADY,
    S_AXI_GP1_BVALID,
    S_AXI_GP1_RLAST,
    S_AXI_GP1_RVALID,
    S_AXI_GP1_WREADY,
    S_AXI_GP1_BRESP,
    S_AXI_GP1_RRESP,
    S_AXI_GP1_RDATA,
    S_AXI_GP1_BID,
    S_AXI_GP1_RID,
    S_AXI_GP1_ACLK,
    S_AXI_GP1_ARVALID,
    S_AXI_GP1_AWVALID,
    S_AXI_GP1_BREADY,
    S_AXI_GP1_RREADY,
    S_AXI_GP1_WLAST,
    S_AXI_GP1_WVALID,
    S_AXI_GP1_ARBURST,
    S_AXI_GP1_ARLOCK,
    S_AXI_GP1_ARSIZE,
    S_AXI_GP1_AWBURST,
    S_AXI_GP1_AWLOCK,
    S_AXI_GP1_AWSIZE,
    S_AXI_GP1_ARPROT,
    S_AXI_GP1_AWPROT,
    S_AXI_GP1_ARADDR,
    S_AXI_GP1_AWADDR,
    S_AXI_GP1_WDATA,
    S_AXI_GP1_ARCACHE,
    S_AXI_GP1_ARLEN,
    S_AXI_GP1_ARQOS,
    S_AXI_GP1_AWCACHE,
    S_AXI_GP1_AWLEN,
    S_AXI_GP1_AWQOS,
    S_AXI_GP1_WSTRB,
    S_AXI_GP1_ARID,
    S_AXI_GP1_AWID,
    S_AXI_GP1_WID,
    S_AXI_ACP_ARESETN,
    S_AXI_ACP_AWREADY,
    S_AXI_ACP_ARREADY,
    S_AXI_ACP_BVALID,
    S_AXI_ACP_RLAST,
    S_AXI_ACP_RVALID,
    S_AXI_ACP_WREADY,
    S_AXI_ACP_BRESP,
    S_AXI_ACP_RRESP,
    S_AXI_ACP_BID,
    S_AXI_ACP_RID,
    S_AXI_ACP_RDATA,
    S_AXI_ACP_ACLK,
    S_AXI_ACP_ARVALID,
    S_AXI_ACP_AWVALID,
    S_AXI_ACP_BREADY,
    S_AXI_ACP_RREADY,
    S_AXI_ACP_WLAST,
    S_AXI_ACP_WVALID,
    S_AXI_ACP_ARID,
    S_AXI_ACP_ARPROT,
    S_AXI_ACP_AWID,
    S_AXI_ACP_AWPROT,
    S_AXI_ACP_WID,
    S_AXI_ACP_ARADDR,
    S_AXI_ACP_AWADDR,
    S_AXI_ACP_ARCACHE,
    S_AXI_ACP_ARLEN,
    S_AXI_ACP_ARQOS,
    S_AXI_ACP_AWCACHE,
    S_AXI_ACP_AWLEN,
    S_AXI_ACP_AWQOS,
    S_AXI_ACP_ARBURST,
    S_AXI_ACP_ARLOCK,
    S_AXI_ACP_ARSIZE,
    S_AXI_ACP_AWBURST,
    S_AXI_ACP_AWLOCK,
    S_AXI_ACP_AWSIZE,
    S_AXI_ACP_ARUSER,
    S_AXI_ACP_AWUSER,
    S_AXI_ACP_WDATA,
    S_AXI_ACP_WSTRB,
    S_AXI_HP0_ARESETN,
    S_AXI_HP0_ARREADY,
    S_AXI_HP0_AWREADY,
    S_AXI_HP0_BVALID,
    S_AXI_HP0_RLAST,
    S_AXI_HP0_RVALID,
    S_AXI_HP0_WREADY,
    S_AXI_HP0_BRESP,
    S_AXI_HP0_RRESP,
    S_AXI_HP0_BID,
    S_AXI_HP0_RID,
    S_AXI_HP0_RDATA,
    S_AXI_HP0_RCOUNT,
    S_AXI_HP0_WCOUNT,
    S_AXI_HP0_RACOUNT,
    S_AXI_HP0_WACOUNT,
    S_AXI_HP0_ACLK,
    S_AXI_HP0_ARVALID,
    S_AXI_HP0_AWVALID,
    S_AXI_HP0_BREADY,
    S_AXI_HP0_RDISSUECAP1_EN,
    S_AXI_HP0_RREADY,
    S_AXI_HP0_WLAST,
    S_AXI_HP0_WRISSUECAP1_EN,
    S_AXI_HP0_WVALID,
    S_AXI_HP0_ARBURST,
    S_AXI_HP0_ARLOCK,
    S_AXI_HP0_ARSIZE,
    S_AXI_HP0_AWBURST,
    S_AXI_HP0_AWLOCK,
    S_AXI_HP0_AWSIZE,
    S_AXI_HP0_ARPROT,
    S_AXI_HP0_AWPROT,
    S_AXI_HP0_ARADDR,
    S_AXI_HP0_AWADDR,
    S_AXI_HP0_ARCACHE,
    S_AXI_HP0_ARLEN,
    S_AXI_HP0_ARQOS,
    S_AXI_HP0_AWCACHE,
    S_AXI_HP0_AWLEN,
    S_AXI_HP0_AWQOS,
    S_AXI_HP0_ARID,
    S_AXI_HP0_AWID,
    S_AXI_HP0_WID,
    S_AXI_HP0_WDATA,
    S_AXI_HP0_WSTRB,
    S_AXI_HP1_ARESETN,
    S_AXI_HP1_ARREADY,
    S_AXI_HP1_AWREADY,
    S_AXI_HP1_BVALID,
    S_AXI_HP1_RLAST,
    S_AXI_HP1_RVALID,
    S_AXI_HP1_WREADY,
    S_AXI_HP1_BRESP,
    S_AXI_HP1_RRESP,
    S_AXI_HP1_BID,
    S_AXI_HP1_RID,
    S_AXI_HP1_RDATA,
    S_AXI_HP1_RCOUNT,
    S_AXI_HP1_WCOUNT,
    S_AXI_HP1_RACOUNT,
    S_AXI_HP1_WACOUNT,
    S_AXI_HP1_ACLK,
    S_AXI_HP1_ARVALID,
    S_AXI_HP1_AWVALID,
    S_AXI_HP1_BREADY,
    S_AXI_HP1_RDISSUECAP1_EN,
    S_AXI_HP1_RREADY,
    S_AXI_HP1_WLAST,
    S_AXI_HP1_WRISSUECAP1_EN,
    S_AXI_HP1_WVALID,
    S_AXI_HP1_ARBURST,
    S_AXI_HP1_ARLOCK,
    S_AXI_HP1_ARSIZE,
    S_AXI_HP1_AWBURST,
    S_AXI_HP1_AWLOCK,
    S_AXI_HP1_AWSIZE,
    S_AXI_HP1_ARPROT,
    S_AXI_HP1_AWPROT,
    S_AXI_HP1_ARADDR,
    S_AXI_HP1_AWADDR,
    S_AXI_HP1_ARCACHE,
    S_AXI_HP1_ARLEN,
    S_AXI_HP1_ARQOS,
    S_AXI_HP1_AWCACHE,
    S_AXI_HP1_AWLEN,
    S_AXI_HP1_AWQOS,
    S_AXI_HP1_ARID,
    S_AXI_HP1_AWID,
    S_AXI_HP1_WID,
    S_AXI_HP1_WDATA,
    S_AXI_HP1_WSTRB,
    S_AXI_HP2_ARESETN,
    S_AXI_HP2_ARREADY,
    S_AXI_HP2_AWREADY,
    S_AXI_HP2_BVALID,
    S_AXI_HP2_RLAST,
    S_AXI_HP2_RVALID,
    S_AXI_HP2_WREADY,
    S_AXI_HP2_BRESP,
    S_AXI_HP2_RRESP,
    S_AXI_HP2_BID,
    S_AXI_HP2_RID,
    S_AXI_HP2_RDATA,
    S_AXI_HP2_RCOUNT,
    S_AXI_HP2_WCOUNT,
    S_AXI_HP2_RACOUNT,
    S_AXI_HP2_WACOUNT,
    S_AXI_HP2_ACLK,
    S_AXI_HP2_ARVALID,
    S_AXI_HP2_AWVALID,
    S_AXI_HP2_BREADY,
    S_AXI_HP2_RDISSUECAP1_EN,
    S_AXI_HP2_RREADY,
    S_AXI_HP2_WLAST,
    S_AXI_HP2_WRISSUECAP1_EN,
    S_AXI_HP2_WVALID,
    S_AXI_HP2_ARBURST,
    S_AXI_HP2_ARLOCK,
    S_AXI_HP2_ARSIZE,
    S_AXI_HP2_AWBURST,
    S_AXI_HP2_AWLOCK,
    S_AXI_HP2_AWSIZE,
    S_AXI_HP2_ARPROT,
    S_AXI_HP2_AWPROT,
    S_AXI_HP2_ARADDR,
    S_AXI_HP2_AWADDR,
    S_AXI_HP2_ARCACHE,
    S_AXI_HP2_ARLEN,
    S_AXI_HP2_ARQOS,
    S_AXI_HP2_AWCACHE,
    S_AXI_HP2_AWLEN,
    S_AXI_HP2_AWQOS,
    S_AXI_HP2_ARID,
    S_AXI_HP2_AWID,
    S_AXI_HP2_WID,
    S_AXI_HP2_WDATA,
    S_AXI_HP2_WSTRB,
    S_AXI_HP3_ARESETN,
    S_AXI_HP3_ARREADY,
    S_AXI_HP3_AWREADY,
    S_AXI_HP3_BVALID,
    S_AXI_HP3_RLAST,
    S_AXI_HP3_RVALID,
    S_AXI_HP3_WREADY,
    S_AXI_HP3_BRESP,
    S_AXI_HP3_RRESP,
    S_AXI_HP3_BID,
    S_AXI_HP3_RID,
    S_AXI_HP3_RDATA,
    S_AXI_HP3_RCOUNT,
    S_AXI_HP3_WCOUNT,
    S_AXI_HP3_RACOUNT,
    S_AXI_HP3_WACOUNT,
    S_AXI_HP3_ACLK,
    S_AXI_HP3_ARVALID,
    S_AXI_HP3_AWVALID,
    S_AXI_HP3_BREADY,
    S_AXI_HP3_RDISSUECAP1_EN,
    S_AXI_HP3_RREADY,
    S_AXI_HP3_WLAST,
    S_AXI_HP3_WRISSUECAP1_EN,
    S_AXI_HP3_WVALID,
    S_AXI_HP3_ARBURST,
    S_AXI_HP3_ARLOCK,
    S_AXI_HP3_ARSIZE,
    S_AXI_HP3_AWBURST,
    S_AXI_HP3_AWLOCK,
    S_AXI_HP3_AWSIZE,
    S_AXI_HP3_ARPROT,
    S_AXI_HP3_AWPROT,
    S_AXI_HP3_ARADDR,
    S_AXI_HP3_AWADDR,
    S_AXI_HP3_ARCACHE,
    S_AXI_HP3_ARLEN,
    S_AXI_HP3_ARQOS,
    S_AXI_HP3_AWCACHE,
    S_AXI_HP3_AWLEN,
    S_AXI_HP3_AWQOS,
    S_AXI_HP3_ARID,
    S_AXI_HP3_AWID,
    S_AXI_HP3_WID,
    S_AXI_HP3_WDATA,
    S_AXI_HP3_WSTRB,
    DMA0_DATYPE,
    DMA0_DAVALID,
    DMA0_DRREADY,
    DMA0_RSTN,
    DMA0_ACLK,
    DMA0_DAREADY,
    DMA0_DRLAST,
    DMA0_DRVALID,
    DMA0_DRTYPE,
    DMA1_DATYPE,
    DMA1_DAVALID,
    DMA1_DRREADY,
    DMA1_RSTN,
    DMA1_ACLK,
    DMA1_DAREADY,
    DMA1_DRLAST,
    DMA1_DRVALID,
    DMA1_DRTYPE,
    DMA2_DATYPE,
    DMA2_DAVALID,
    DMA2_DRREADY,
    DMA2_RSTN,
    DMA2_ACLK,
    DMA2_DAREADY,
    DMA2_DRLAST,
    DMA2_DRVALID,
    DMA3_DRVALID,
    DMA3_DATYPE,
    DMA3_DAVALID,
    DMA3_DRREADY,
    DMA3_RSTN,
    DMA3_ACLK,
    DMA3_DAREADY,
    DMA3_DRLAST,
    DMA2_DRTYPE,
    DMA3_DRTYPE,
    FTMD_TRACEIN_DATA,
    FTMD_TRACEIN_VALID,
    FTMD_TRACEIN_CLK,
    FTMD_TRACEIN_ATID,
    FTMT_F2P_TRIG,
    FTMT_F2P_TRIGACK,
    FTMT_F2P_DEBUG,
    FTMT_P2F_TRIGACK,
    FTMT_P2F_TRIG,
    FTMT_P2F_DEBUG,
    FCLK_CLK3,
    FCLK_CLK2,
    FCLK_CLK1,
    FCLK_CLK0,
    FCLK_CLKTRIG3_N,
    FCLK_CLKTRIG2_N,
    FCLK_CLKTRIG1_N,
    FCLK_CLKTRIG0_N,
    FCLK_RESET3_N,
    FCLK_RESET2_N,
    FCLK_RESET1_N,
    FCLK_RESET0_N,
    FPGA_IDLE_N,
    DDR_ARB,
    IRQ_F2P,
    Core0_nFIQ,
    Core0_nIRQ,
    Core1_nFIQ,
    Core1_nIRQ,
    EVENT_EVENTO,
    EVENT_STANDBYWFE,
    EVENT_STANDBYWFI,
    EVENT_EVENTI,
    MIO,
    DDR_Clk,
    DDR_Clk_n,
    DDR_CKE,
    DDR_CS_n,
    DDR_RAS_n,
    DDR_CAS_n,
    DDR_WEB,
    DDR_BankAddr,
    DDR_Addr,
    DDR_ODT,
    DDR_DRSTB,
    DDR_DQ,
    DDR_DM,
    DDR_DQS,
    DDR_DQS_n,
    DDR_VRN,
    DDR_VRP,
    PS_SRSTB,
    PS_CLK,
    PS_PORB,
    IRQ_P2F_DMAC_ABORT,
    IRQ_P2F_DMAC0,
    IRQ_P2F_DMAC1,
    IRQ_P2F_DMAC2,
    IRQ_P2F_DMAC3,
    IRQ_P2F_DMAC4,
    IRQ_P2F_DMAC5,
    IRQ_P2F_DMAC6,
    IRQ_P2F_DMAC7,
    IRQ_P2F_SMC,
    IRQ_P2F_QSPI,
    IRQ_P2F_CTI,
    IRQ_P2F_GPIO,
    IRQ_P2F_USB0,
    IRQ_P2F_ENET0,
    IRQ_P2F_ENET_WAKE0,
    IRQ_P2F_SDIO0,
    IRQ_P2F_I2C0,
    IRQ_P2F_SPI0,
    IRQ_P2F_UART0,
    IRQ_P2F_CAN0,
    IRQ_P2F_USB1,
    IRQ_P2F_ENET1,
    IRQ_P2F_ENET_WAKE1,
    IRQ_P2F_SDIO1,
    IRQ_P2F_I2C1,
    IRQ_P2F_SPI1,
    IRQ_P2F_UART1,
    IRQ_P2F_CAN1
  );
  output CAN0_PHY_TX;
  input CAN0_PHY_RX;
  output CAN1_PHY_TX;
  input CAN1_PHY_RX;
  output ENET0_GMII_TX_EN;
  output ENET0_GMII_TX_ER;
  output ENET0_MDIO_MDC;
  output ENET0_MDIO_O;
  output ENET0_MDIO_T;
  output ENET0_PTP_DELAY_REQ_RX;
  output ENET0_PTP_DELAY_REQ_TX;
  output ENET0_PTP_PDELAY_REQ_RX;
  output ENET0_PTP_PDELAY_REQ_TX;
  output ENET0_PTP_PDELAY_RESP_RX;
  output ENET0_PTP_PDELAY_RESP_TX;
  output ENET0_PTP_SYNC_FRAME_RX;
  output ENET0_PTP_SYNC_FRAME_TX;
  output ENET0_SOF_RX;
  output ENET0_SOF_TX;
  output [7:0] ENET0_GMII_TXD;
  input ENET0_GMII_COL;
  input ENET0_GMII_CRS;
  input ENET0_EXT_INTIN;
  input ENET0_GMII_RX_CLK;
  input ENET0_GMII_RX_DV;
  input ENET0_GMII_RX_ER;
  input ENET0_GMII_TX_CLK;
  input ENET0_MDIO_I;
  input [7:0] ENET0_GMII_RXD;
  output ENET1_GMII_TX_EN;
  output ENET1_GMII_TX_ER;
  output ENET1_MDIO_MDC;
  output ENET1_MDIO_O;
  output ENET1_MDIO_T;
  output ENET1_PTP_DELAY_REQ_RX;
  output ENET1_PTP_DELAY_REQ_TX;
  output ENET1_PTP_PDELAY_REQ_RX;
  output ENET1_PTP_PDELAY_REQ_TX;
  output ENET1_PTP_PDELAY_RESP_RX;
  output ENET1_PTP_PDELAY_RESP_TX;
  output ENET1_PTP_SYNC_FRAME_RX;
  output ENET1_PTP_SYNC_FRAME_TX;
  output ENET1_SOF_RX;
  output ENET1_SOF_TX;
  output [7:0] ENET1_GMII_TXD;
  input ENET1_GMII_COL;
  input ENET1_GMII_CRS;
  input ENET1_EXT_INTIN;
  input ENET1_GMII_RX_CLK;
  input ENET1_GMII_RX_DV;
  input ENET1_GMII_RX_ER;
  input ENET1_GMII_TX_CLK;
  input ENET1_MDIO_I;
  input [7:0] ENET1_GMII_RXD;
  input [63:0] GPIO_I;
  output [63:0] GPIO_O;
  output [63:0] GPIO_T;
  input I2C0_SDA_I;
  output I2C0_SDA_O;
  output I2C0_SDA_T;
  input I2C0_SCL_I;
  output I2C0_SCL_O;
  output I2C0_SCL_T;
  input I2C1_SDA_I;
  output I2C1_SDA_O;
  output I2C1_SDA_T;
  input I2C1_SCL_I;
  output I2C1_SCL_O;
  output I2C1_SCL_T;
  input PJTAG_TCK;
  input PJTAG_TMS;
  input PJTAG_TD_I;
  output PJTAG_TD_T;
  output PJTAG_TD_O;
  output SDIO0_CLK;
  input SDIO0_CLK_FB;
  output SDIO0_CMD_O;
  input SDIO0_CMD_I;
  output SDIO0_CMD_T;
  input [3:0] SDIO0_DATA_I;
  output [3:0] SDIO0_DATA_O;
  output [3:0] SDIO0_DATA_T;
  output SDIO0_LED;
  input SDIO0_CDN;
  input SDIO0_WP;
  output SDIO0_BUSPOW;
  output [2:0] SDIO0_BUSVOLT;
  output SDIO1_CLK;
  input SDIO1_CLK_FB;
  output SDIO1_CMD_O;
  input SDIO1_CMD_I;
  output SDIO1_CMD_T;
  input [3:0] SDIO1_DATA_I;
  output [3:0] SDIO1_DATA_O;
  output [3:0] SDIO1_DATA_T;
  output SDIO1_LED;
  input SDIO1_CDN;
  input SDIO1_WP;
  output SDIO1_BUSPOW;
  output [2:0] SDIO1_BUSVOLT;
  input SPI0_SCLK_I;
  output SPI0_SCLK_O;
  output SPI0_SCLK_T;
  input SPI0_MOSI_I;
  output SPI0_MOSI_O;
  output SPI0_MOSI_T;
  input SPI0_MISO_I;
  output SPI0_MISO_O;
  output SPI0_MISO_T;
  input SPI0_SS_I;
  output SPI0_SS_O;
  output SPI0_SS1_O;
  output SPI0_SS2_O;
  output SPI0_SS_T;
  input SPI1_SCLK_I;
  output SPI1_SCLK_O;
  output SPI1_SCLK_T;
  input SPI1_MOSI_I;
  output SPI1_MOSI_O;
  output SPI1_MOSI_T;
  input SPI1_MISO_I;
  output SPI1_MISO_O;
  output SPI1_MISO_T;
  input SPI1_SS_I;
  output SPI1_SS_O;
  output SPI1_SS1_O;
  output SPI1_SS2_O;
  output SPI1_SS_T;
  output UART0_DTRN;
  output UART0_RTSN;
  output UART0_TX;
  input UART0_CTSN;
  input UART0_DCDN;
  input UART0_DSRN;
  input UART0_RIN;
  input UART0_RX;
  output UART1_DTRN;
  output UART1_RTSN;
  output UART1_TX;
  input UART1_CTSN;
  input UART1_DCDN;
  input UART1_DSRN;
  input UART1_RIN;
  input UART1_RX;
  output TTC0_WAVE0_OUT;
  output TTC0_WAVE1_OUT;
  output TTC0_WAVE2_OUT;
  input TTC0_CLK0_IN;
  input TTC0_CLK1_IN;
  input TTC0_CLK2_IN;
  output TTC1_WAVE0_OUT;
  output TTC1_WAVE1_OUT;
  output TTC1_WAVE2_OUT;
  input TTC1_CLK0_IN;
  input TTC1_CLK1_IN;
  input TTC1_CLK2_IN;
  input WDT_CLK_IN;
  output WDT_RST_OUT;
  input TRACE_CLK;
  output TRACE_CTL;
  output [31:0] TRACE_DATA;
  output [1:0] USB0_PORT_INDCTL;
  output [1:0] USB1_PORT_INDCTL;
  output USB0_VBUS_PWRSELECT;
  output USB1_VBUS_PWRSELECT;
  input USB0_VBUS_PWRFAULT;
  input USB1_VBUS_PWRFAULT;
  input SRAM_INTIN;
  output M_AXI_GP0_ARESETN;
  output M_AXI_GP0_ARVALID;
  output M_AXI_GP0_AWVALID;
  output M_AXI_GP0_BREADY;
  output M_AXI_GP0_RREADY;
  output M_AXI_GP0_WLAST;
  output M_AXI_GP0_WVALID;
  output [11:0] M_AXI_GP0_ARID;
  output [11:0] M_AXI_GP0_AWID;
  output [11:0] M_AXI_GP0_WID;
  output [1:0] M_AXI_GP0_ARBURST;
  output [1:0] M_AXI_GP0_ARLOCK;
  output [2:0] M_AXI_GP0_ARSIZE;
  output [1:0] M_AXI_GP0_AWBURST;
  output [1:0] M_AXI_GP0_AWLOCK;
  output [2:0] M_AXI_GP0_AWSIZE;
  output [2:0] M_AXI_GP0_ARPROT;
  output [2:0] M_AXI_GP0_AWPROT;
  output [31:0] M_AXI_GP0_ARADDR;
  output [31:0] M_AXI_GP0_AWADDR;
  output [31:0] M_AXI_GP0_WDATA;
  output [3:0] M_AXI_GP0_ARCACHE;
  output [3:0] M_AXI_GP0_ARLEN;
  output [3:0] M_AXI_GP0_ARQOS;
  output [3:0] M_AXI_GP0_AWCACHE;
  output [3:0] M_AXI_GP0_AWLEN;
  output [3:0] M_AXI_GP0_AWQOS;
  output [3:0] M_AXI_GP0_WSTRB;
  input M_AXI_GP0_ACLK;
  input M_AXI_GP0_ARREADY;
  input M_AXI_GP0_AWREADY;
  input M_AXI_GP0_BVALID;
  input M_AXI_GP0_RLAST;
  input M_AXI_GP0_RVALID;
  input M_AXI_GP0_WREADY;
  input [11:0] M_AXI_GP0_BID;
  input [11:0] M_AXI_GP0_RID;
  input [1:0] M_AXI_GP0_BRESP;
  input [1:0] M_AXI_GP0_RRESP;
  input [31:0] M_AXI_GP0_RDATA;
  output M_AXI_GP1_ARESETN;
  output M_AXI_GP1_ARVALID;
  output M_AXI_GP1_AWVALID;
  output M_AXI_GP1_BREADY;
  output M_AXI_GP1_RREADY;
  output M_AXI_GP1_WLAST;
  output M_AXI_GP1_WVALID;
  output [11:0] M_AXI_GP1_ARID;
  output [11:0] M_AXI_GP1_AWID;
  output [11:0] M_AXI_GP1_WID;
  output [1:0] M_AXI_GP1_ARBURST;
  output [1:0] M_AXI_GP1_ARLOCK;
  output [2:0] M_AXI_GP1_ARSIZE;
  output [1:0] M_AXI_GP1_AWBURST;
  output [1:0] M_AXI_GP1_AWLOCK;
  output [2:0] M_AXI_GP1_AWSIZE;
  output [2:0] M_AXI_GP1_ARPROT;
  output [2:0] M_AXI_GP1_AWPROT;
  output [31:0] M_AXI_GP1_ARADDR;
  output [31:0] M_AXI_GP1_AWADDR;
  output [31:0] M_AXI_GP1_WDATA;
  output [3:0] M_AXI_GP1_ARCACHE;
  output [3:0] M_AXI_GP1_ARLEN;
  output [3:0] M_AXI_GP1_ARQOS;
  output [3:0] M_AXI_GP1_AWCACHE;
  output [3:0] M_AXI_GP1_AWLEN;
  output [3:0] M_AXI_GP1_AWQOS;
  output [3:0] M_AXI_GP1_WSTRB;
  input M_AXI_GP1_ACLK;
  input M_AXI_GP1_ARREADY;
  input M_AXI_GP1_AWREADY;
  input M_AXI_GP1_BVALID;
  input M_AXI_GP1_RLAST;
  input M_AXI_GP1_RVALID;
  input M_AXI_GP1_WREADY;
  input [11:0] M_AXI_GP1_BID;
  input [11:0] M_AXI_GP1_RID;
  input [1:0] M_AXI_GP1_BRESP;
  input [1:0] M_AXI_GP1_RRESP;
  input [31:0] M_AXI_GP1_RDATA;
  output S_AXI_GP0_ARESETN;
  output S_AXI_GP0_ARREADY;
  output S_AXI_GP0_AWREADY;
  output S_AXI_GP0_BVALID;
  output S_AXI_GP0_RLAST;
  output S_AXI_GP0_RVALID;
  output S_AXI_GP0_WREADY;
  output [1:0] S_AXI_GP0_BRESP;
  output [1:0] S_AXI_GP0_RRESP;
  output [31:0] S_AXI_GP0_RDATA;
  output [5:0] S_AXI_GP0_BID;
  output [5:0] S_AXI_GP0_RID;
  input S_AXI_GP0_ACLK;
  input S_AXI_GP0_ARVALID;
  input S_AXI_GP0_AWVALID;
  input S_AXI_GP0_BREADY;
  input S_AXI_GP0_RREADY;
  input S_AXI_GP0_WLAST;
  input S_AXI_GP0_WVALID;
  input [1:0] S_AXI_GP0_ARBURST;
  input [1:0] S_AXI_GP0_ARLOCK;
  input [2:0] S_AXI_GP0_ARSIZE;
  input [1:0] S_AXI_GP0_AWBURST;
  input [1:0] S_AXI_GP0_AWLOCK;
  input [2:0] S_AXI_GP0_AWSIZE;
  input [2:0] S_AXI_GP0_ARPROT;
  input [2:0] S_AXI_GP0_AWPROT;
  input [31:0] S_AXI_GP0_ARADDR;
  input [31:0] S_AXI_GP0_AWADDR;
  input [31:0] S_AXI_GP0_WDATA;
  input [3:0] S_AXI_GP0_ARCACHE;
  input [3:0] S_AXI_GP0_ARLEN;
  input [3:0] S_AXI_GP0_ARQOS;
  input [3:0] S_AXI_GP0_AWCACHE;
  input [3:0] S_AXI_GP0_AWLEN;
  input [3:0] S_AXI_GP0_AWQOS;
  input [3:0] S_AXI_GP0_WSTRB;
  input [5:0] S_AXI_GP0_ARID;
  input [5:0] S_AXI_GP0_AWID;
  input [5:0] S_AXI_GP0_WID;
  output S_AXI_GP1_ARESETN;
  output S_AXI_GP1_ARREADY;
  output S_AXI_GP1_AWREADY;
  output S_AXI_GP1_BVALID;
  output S_AXI_GP1_RLAST;
  output S_AXI_GP1_RVALID;
  output S_AXI_GP1_WREADY;
  output [1:0] S_AXI_GP1_BRESP;
  output [1:0] S_AXI_GP1_RRESP;
  output [31:0] S_AXI_GP1_RDATA;
  output [5:0] S_AXI_GP1_BID;
  output [5:0] S_AXI_GP1_RID;
  input S_AXI_GP1_ACLK;
  input S_AXI_GP1_ARVALID;
  input S_AXI_GP1_AWVALID;
  input S_AXI_GP1_BREADY;
  input S_AXI_GP1_RREADY;
  input S_AXI_GP1_WLAST;
  input S_AXI_GP1_WVALID;
  input [1:0] S_AXI_GP1_ARBURST;
  input [1:0] S_AXI_GP1_ARLOCK;
  input [2:0] S_AXI_GP1_ARSIZE;
  input [1:0] S_AXI_GP1_AWBURST;
  input [1:0] S_AXI_GP1_AWLOCK;
  input [2:0] S_AXI_GP1_AWSIZE;
  input [2:0] S_AXI_GP1_ARPROT;
  input [2:0] S_AXI_GP1_AWPROT;
  input [31:0] S_AXI_GP1_ARADDR;
  input [31:0] S_AXI_GP1_AWADDR;
  input [31:0] S_AXI_GP1_WDATA;
  input [3:0] S_AXI_GP1_ARCACHE;
  input [3:0] S_AXI_GP1_ARLEN;
  input [3:0] S_AXI_GP1_ARQOS;
  input [3:0] S_AXI_GP1_AWCACHE;
  input [3:0] S_AXI_GP1_AWLEN;
  input [3:0] S_AXI_GP1_AWQOS;
  input [3:0] S_AXI_GP1_WSTRB;
  input [5:0] S_AXI_GP1_ARID;
  input [5:0] S_AXI_GP1_AWID;
  input [5:0] S_AXI_GP1_WID;
  output S_AXI_ACP_ARESETN;
  output S_AXI_ACP_AWREADY;
  output S_AXI_ACP_ARREADY;
  output S_AXI_ACP_BVALID;
  output S_AXI_ACP_RLAST;
  output S_AXI_ACP_RVALID;
  output S_AXI_ACP_WREADY;
  output [1:0] S_AXI_ACP_BRESP;
  output [1:0] S_AXI_ACP_RRESP;
  output [2:0] S_AXI_ACP_BID;
  output [2:0] S_AXI_ACP_RID;
  output [63:0] S_AXI_ACP_RDATA;
  input S_AXI_ACP_ACLK;
  input S_AXI_ACP_ARVALID;
  input S_AXI_ACP_AWVALID;
  input S_AXI_ACP_BREADY;
  input S_AXI_ACP_RREADY;
  input S_AXI_ACP_WLAST;
  input S_AXI_ACP_WVALID;
  input [2:0] S_AXI_ACP_ARID;
  input [2:0] S_AXI_ACP_ARPROT;
  input [2:0] S_AXI_ACP_AWID;
  input [2:0] S_AXI_ACP_AWPROT;
  input [2:0] S_AXI_ACP_WID;
  input [31:0] S_AXI_ACP_ARADDR;
  input [31:0] S_AXI_ACP_AWADDR;
  input [3:0] S_AXI_ACP_ARCACHE;
  input [3:0] S_AXI_ACP_ARLEN;
  input [3:0] S_AXI_ACP_ARQOS;
  input [3:0] S_AXI_ACP_AWCACHE;
  input [3:0] S_AXI_ACP_AWLEN;
  input [3:0] S_AXI_ACP_AWQOS;
  input [1:0] S_AXI_ACP_ARBURST;
  input [1:0] S_AXI_ACP_ARLOCK;
  input [2:0] S_AXI_ACP_ARSIZE;
  input [1:0] S_AXI_ACP_AWBURST;
  input [1:0] S_AXI_ACP_AWLOCK;
  input [2:0] S_AXI_ACP_AWSIZE;
  input [4:0] S_AXI_ACP_ARUSER;
  input [4:0] S_AXI_ACP_AWUSER;
  input [63:0] S_AXI_ACP_WDATA;
  input [7:0] S_AXI_ACP_WSTRB;
  output S_AXI_HP0_ARESETN;
  output S_AXI_HP0_ARREADY;
  output S_AXI_HP0_AWREADY;
  output S_AXI_HP0_BVALID;
  output S_AXI_HP0_RLAST;
  output S_AXI_HP0_RVALID;
  output S_AXI_HP0_WREADY;
  output [1:0] S_AXI_HP0_BRESP;
  output [1:0] S_AXI_HP0_RRESP;
  output [1:0] S_AXI_HP0_BID;
  output [1:0] S_AXI_HP0_RID;
  output [63:0] S_AXI_HP0_RDATA;
  output [7:0] S_AXI_HP0_RCOUNT;
  output [7:0] S_AXI_HP0_WCOUNT;
  output [2:0] S_AXI_HP0_RACOUNT;
  output [5:0] S_AXI_HP0_WACOUNT;
  input S_AXI_HP0_ACLK;
  input S_AXI_HP0_ARVALID;
  input S_AXI_HP0_AWVALID;
  input S_AXI_HP0_BREADY;
  input S_AXI_HP0_RDISSUECAP1_EN;
  input S_AXI_HP0_RREADY;
  input S_AXI_HP0_WLAST;
  input S_AXI_HP0_WRISSUECAP1_EN;
  input S_AXI_HP0_WVALID;
  input [1:0] S_AXI_HP0_ARBURST;
  input [1:0] S_AXI_HP0_ARLOCK;
  input [2:0] S_AXI_HP0_ARSIZE;
  input [1:0] S_AXI_HP0_AWBURST;
  input [1:0] S_AXI_HP0_AWLOCK;
  input [2:0] S_AXI_HP0_AWSIZE;
  input [2:0] S_AXI_HP0_ARPROT;
  input [2:0] S_AXI_HP0_AWPROT;
  input [31:0] S_AXI_HP0_ARADDR;
  input [31:0] S_AXI_HP0_AWADDR;
  input [3:0] S_AXI_HP0_ARCACHE;
  input [3:0] S_AXI_HP0_ARLEN;
  input [3:0] S_AXI_HP0_ARQOS;
  input [3:0] S_AXI_HP0_AWCACHE;
  input [3:0] S_AXI_HP0_AWLEN;
  input [3:0] S_AXI_HP0_AWQOS;
  input [1:0] S_AXI_HP0_ARID;
  input [1:0] S_AXI_HP0_AWID;
  input [1:0] S_AXI_HP0_WID;
  input [63:0] S_AXI_HP0_WDATA;
  input [7:0] S_AXI_HP0_WSTRB;
  output S_AXI_HP1_ARESETN;
  output S_AXI_HP1_ARREADY;
  output S_AXI_HP1_AWREADY;
  output S_AXI_HP1_BVALID;
  output S_AXI_HP1_RLAST;
  output S_AXI_HP1_RVALID;
  output S_AXI_HP1_WREADY;
  output [1:0] S_AXI_HP1_BRESP;
  output [1:0] S_AXI_HP1_RRESP;
  output [5:0] S_AXI_HP1_BID;
  output [5:0] S_AXI_HP1_RID;
  output [63:0] S_AXI_HP1_RDATA;
  output [7:0] S_AXI_HP1_RCOUNT;
  output [7:0] S_AXI_HP1_WCOUNT;
  output [2:0] S_AXI_HP1_RACOUNT;
  output [5:0] S_AXI_HP1_WACOUNT;
  input S_AXI_HP1_ACLK;
  input S_AXI_HP1_ARVALID;
  input S_AXI_HP1_AWVALID;
  input S_AXI_HP1_BREADY;
  input S_AXI_HP1_RDISSUECAP1_EN;
  input S_AXI_HP1_RREADY;
  input S_AXI_HP1_WLAST;
  input S_AXI_HP1_WRISSUECAP1_EN;
  input S_AXI_HP1_WVALID;
  input [1:0] S_AXI_HP1_ARBURST;
  input [1:0] S_AXI_HP1_ARLOCK;
  input [2:0] S_AXI_HP1_ARSIZE;
  input [1:0] S_AXI_HP1_AWBURST;
  input [1:0] S_AXI_HP1_AWLOCK;
  input [2:0] S_AXI_HP1_AWSIZE;
  input [2:0] S_AXI_HP1_ARPROT;
  input [2:0] S_AXI_HP1_AWPROT;
  input [31:0] S_AXI_HP1_ARADDR;
  input [31:0] S_AXI_HP1_AWADDR;
  input [3:0] S_AXI_HP1_ARCACHE;
  input [3:0] S_AXI_HP1_ARLEN;
  input [3:0] S_AXI_HP1_ARQOS;
  input [3:0] S_AXI_HP1_AWCACHE;
  input [3:0] S_AXI_HP1_AWLEN;
  input [3:0] S_AXI_HP1_AWQOS;
  input [5:0] S_AXI_HP1_ARID;
  input [5:0] S_AXI_HP1_AWID;
  input [5:0] S_AXI_HP1_WID;
  input [63:0] S_AXI_HP1_WDATA;
  input [7:0] S_AXI_HP1_WSTRB;
  output S_AXI_HP2_ARESETN;
  output S_AXI_HP2_ARREADY;
  output S_AXI_HP2_AWREADY;
  output S_AXI_HP2_BVALID;
  output S_AXI_HP2_RLAST;
  output S_AXI_HP2_RVALID;
  output S_AXI_HP2_WREADY;
  output [1:0] S_AXI_HP2_BRESP;
  output [1:0] S_AXI_HP2_RRESP;
  output [5:0] S_AXI_HP2_BID;
  output [5:0] S_AXI_HP2_RID;
  output [63:0] S_AXI_HP2_RDATA;
  output [7:0] S_AXI_HP2_RCOUNT;
  output [7:0] S_AXI_HP2_WCOUNT;
  output [2:0] S_AXI_HP2_RACOUNT;
  output [5:0] S_AXI_HP2_WACOUNT;
  input S_AXI_HP2_ACLK;
  input S_AXI_HP2_ARVALID;
  input S_AXI_HP2_AWVALID;
  input S_AXI_HP2_BREADY;
  input S_AXI_HP2_RDISSUECAP1_EN;
  input S_AXI_HP2_RREADY;
  input S_AXI_HP2_WLAST;
  input S_AXI_HP2_WRISSUECAP1_EN;
  input S_AXI_HP2_WVALID;
  input [1:0] S_AXI_HP2_ARBURST;
  input [1:0] S_AXI_HP2_ARLOCK;
  input [2:0] S_AXI_HP2_ARSIZE;
  input [1:0] S_AXI_HP2_AWBURST;
  input [1:0] S_AXI_HP2_AWLOCK;
  input [2:0] S_AXI_HP2_AWSIZE;
  input [2:0] S_AXI_HP2_ARPROT;
  input [2:0] S_AXI_HP2_AWPROT;
  input [31:0] S_AXI_HP2_ARADDR;
  input [31:0] S_AXI_HP2_AWADDR;
  input [3:0] S_AXI_HP2_ARCACHE;
  input [3:0] S_AXI_HP2_ARLEN;
  input [3:0] S_AXI_HP2_ARQOS;
  input [3:0] S_AXI_HP2_AWCACHE;
  input [3:0] S_AXI_HP2_AWLEN;
  input [3:0] S_AXI_HP2_AWQOS;
  input [5:0] S_AXI_HP2_ARID;
  input [5:0] S_AXI_HP2_AWID;
  input [5:0] S_AXI_HP2_WID;
  input [63:0] S_AXI_HP2_WDATA;
  input [7:0] S_AXI_HP2_WSTRB;
  output S_AXI_HP3_ARESETN;
  output S_AXI_HP3_ARREADY;
  output S_AXI_HP3_AWREADY;
  output S_AXI_HP3_BVALID;
  output S_AXI_HP3_RLAST;
  output S_AXI_HP3_RVALID;
  output S_AXI_HP3_WREADY;
  output [1:0] S_AXI_HP3_BRESP;
  output [1:0] S_AXI_HP3_RRESP;
  output [5:0] S_AXI_HP3_BID;
  output [5:0] S_AXI_HP3_RID;
  output [63:0] S_AXI_HP3_RDATA;
  output [7:0] S_AXI_HP3_RCOUNT;
  output [7:0] S_AXI_HP3_WCOUNT;
  output [2:0] S_AXI_HP3_RACOUNT;
  output [5:0] S_AXI_HP3_WACOUNT;
  input S_AXI_HP3_ACLK;
  input S_AXI_HP3_ARVALID;
  input S_AXI_HP3_AWVALID;
  input S_AXI_HP3_BREADY;
  input S_AXI_HP3_RDISSUECAP1_EN;
  input S_AXI_HP3_RREADY;
  input S_AXI_HP3_WLAST;
  input S_AXI_HP3_WRISSUECAP1_EN;
  input S_AXI_HP3_WVALID;
  input [1:0] S_AXI_HP3_ARBURST;
  input [1:0] S_AXI_HP3_ARLOCK;
  input [2:0] S_AXI_HP3_ARSIZE;
  input [1:0] S_AXI_HP3_AWBURST;
  input [1:0] S_AXI_HP3_AWLOCK;
  input [2:0] S_AXI_HP3_AWSIZE;
  input [2:0] S_AXI_HP3_ARPROT;
  input [2:0] S_AXI_HP3_AWPROT;
  input [31:0] S_AXI_HP3_ARADDR;
  input [31:0] S_AXI_HP3_AWADDR;
  input [3:0] S_AXI_HP3_ARCACHE;
  input [3:0] S_AXI_HP3_ARLEN;
  input [3:0] S_AXI_HP3_ARQOS;
  input [3:0] S_AXI_HP3_AWCACHE;
  input [3:0] S_AXI_HP3_AWLEN;
  input [3:0] S_AXI_HP3_AWQOS;
  input [5:0] S_AXI_HP3_ARID;
  input [5:0] S_AXI_HP3_AWID;
  input [5:0] S_AXI_HP3_WID;
  input [63:0] S_AXI_HP3_WDATA;
  input [7:0] S_AXI_HP3_WSTRB;
  output [1:0] DMA0_DATYPE;
  output DMA0_DAVALID;
  output DMA0_DRREADY;
  output DMA0_RSTN;
  input DMA0_ACLK;
  input DMA0_DAREADY;
  input DMA0_DRLAST;
  input DMA0_DRVALID;
  input [1:0] DMA0_DRTYPE;
  output [1:0] DMA1_DATYPE;
  output DMA1_DAVALID;
  output DMA1_DRREADY;
  output DMA1_RSTN;
  input DMA1_ACLK;
  input DMA1_DAREADY;
  input DMA1_DRLAST;
  input DMA1_DRVALID;
  input [1:0] DMA1_DRTYPE;
  output [1:0] DMA2_DATYPE;
  output DMA2_DAVALID;
  output DMA2_DRREADY;
  output DMA2_RSTN;
  input DMA2_ACLK;
  input DMA2_DAREADY;
  input DMA2_DRLAST;
  input DMA2_DRVALID;
  input DMA3_DRVALID;
  output [1:0] DMA3_DATYPE;
  output DMA3_DAVALID;
  output DMA3_DRREADY;
  output DMA3_RSTN;
  input DMA3_ACLK;
  input DMA3_DAREADY;
  input DMA3_DRLAST;
  input [1:0] DMA2_DRTYPE;
  input [1:0] DMA3_DRTYPE;
  input [31:0] FTMD_TRACEIN_DATA;
  input FTMD_TRACEIN_VALID;
  input FTMD_TRACEIN_CLK;
  input [3:0] FTMD_TRACEIN_ATID;
  input [3:0] FTMT_F2P_TRIG;
  output [3:0] FTMT_F2P_TRIGACK;
  input [31:0] FTMT_F2P_DEBUG;
  input [3:0] FTMT_P2F_TRIGACK;
  output [3:0] FTMT_P2F_TRIG;
  output [31:0] FTMT_P2F_DEBUG;
  output FCLK_CLK3;
  output FCLK_CLK2;
  output FCLK_CLK1;
  output FCLK_CLK0;
  input FCLK_CLKTRIG3_N;
  input FCLK_CLKTRIG2_N;
  input FCLK_CLKTRIG1_N;
  input FCLK_CLKTRIG0_N;
  output FCLK_RESET3_N;
  output FCLK_RESET2_N;
  output FCLK_RESET1_N;
  output FCLK_RESET0_N;
  input FPGA_IDLE_N;
  input [3:0] DDR_ARB;
  input [0:0] IRQ_F2P;
  input Core0_nFIQ;
  input Core0_nIRQ;
  input Core1_nFIQ;
  input Core1_nIRQ;
  output EVENT_EVENTO;
  output [1:0] EVENT_STANDBYWFE;
  output [1:0] EVENT_STANDBYWFI;
  input EVENT_EVENTI;
  inout [53:0] MIO;
  inout DDR_Clk;
  inout DDR_Clk_n;
  inout DDR_CKE;
  inout DDR_CS_n;
  inout DDR_RAS_n;
  inout DDR_CAS_n;
  output DDR_WEB;
  inout [2:0] DDR_BankAddr;
  inout [14:0] DDR_Addr;
  inout DDR_ODT;
  inout DDR_DRSTB;
  inout [31:0] DDR_DQ;
  inout [3:0] DDR_DM;
  inout [3:0] DDR_DQS;
  inout [3:0] DDR_DQS_n;
  inout DDR_VRN;
  inout DDR_VRP;
  input PS_SRSTB;
  input PS_CLK;
  input PS_PORB;
  output IRQ_P2F_DMAC_ABORT;
  output IRQ_P2F_DMAC0;
  output IRQ_P2F_DMAC1;
  output IRQ_P2F_DMAC2;
  output IRQ_P2F_DMAC3;
  output IRQ_P2F_DMAC4;
  output IRQ_P2F_DMAC5;
  output IRQ_P2F_DMAC6;
  output IRQ_P2F_DMAC7;
  output IRQ_P2F_SMC;
  output IRQ_P2F_QSPI;
  output IRQ_P2F_CTI;
  output IRQ_P2F_GPIO;
  output IRQ_P2F_USB0;
  output IRQ_P2F_ENET0;
  output IRQ_P2F_ENET_WAKE0;
  output IRQ_P2F_SDIO0;
  output IRQ_P2F_I2C0;
  output IRQ_P2F_SPI0;
  output IRQ_P2F_UART0;
  output IRQ_P2F_CAN0;
  output IRQ_P2F_USB1;
  output IRQ_P2F_ENET1;
  output IRQ_P2F_ENET_WAKE1;
  output IRQ_P2F_SDIO1;
  output IRQ_P2F_I2C1;
  output IRQ_P2F_SPI1;
  output IRQ_P2F_UART1;
  output IRQ_P2F_CAN1;

  (* CORE_GENERATION_INFO = "processing_system7_0,processing_system7,{C_ENET0_PERIPHERAL_ENABLE = 1,C_USB0_PERIPHERAL_ENABLE = 1,C_QSPI_PERIPHERAL_ENABLE = 1,C_DDR_V4.00.A_C_S_AXI_HP3_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP2_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP1_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP0_BASEADDR = 0x00000000,C_DDR_V4.00.A_C_S_AXI_HP3_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP2_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP1_HIGHADDR = 0x3FFFFFFF,C_DDR_V4.00.A_C_S_AXI_HP0_HIGHADDR = 0x3FFFFFFF,C_GPIO_PERIPHERAL_ENABLE = 1,C_GPIO_V2.00.A_C_EN_EMIO_GPIO = 0,C:GPIO_EMIO_GPIO_WIDTH = 64,C_CAN_PERIPHERAL_FREQMHZ = 100,C_FPGA3_PERIPHERAL_FREQMHZ = 25.000000,C_FPGA0_PERIPHERAL_FREQMHZ = 100.000000,C_PRESET_GLOBAL_DEFAULT = powerup,C_FPGA1_PERIPHERAL_FREQMHZ = 150.000000,C_PRESET_GLOBAL_CONFIG = Default,C_PRESET_FPGA_SPEED = -1,C_PRESET_FPGA_PARTNUMBER = xc7z020clg484-1,C_SD0_PERIPHERAL_ENABLE = 1,C_UART1_PERIPHERAL_ENABLE = 1}" *)

  processing_system7
    #(
      .C_EN_EMIO_ENET0 ( 1 ),
      .C_EN_EMIO_ENET1 ( 0 ),
      .C_EN_EMIO_TRACE ( 0 ),
      .C_INCLUDE_TRACE_BUFFER ( 0 ),
      .C_TRACE_BUFFER_FIFO_SIZE ( 128 ),
      .USE_TRACE_DATA_EDGE_DETECTOR ( 0 ),
      .C_TRACE_BUFFER_CLOCK_DELAY ( 12 ),
      .C_EMIO_GPIO_WIDTH ( 64 ),
      .C_INCLUDE_ACP_TRANS_CHECK ( 0 ),
      .C_USE_DEFAULT_ACP_USER_VAL ( 0 ),
      .C_S_AXI_ACP_ARUSER_VAL ( 31 ),
      .C_S_AXI_ACP_AWUSER_VAL ( 31 ),
      .C_DQ_WIDTH ( 32 ),
      .C_DQS_WIDTH ( 4 ),
      .C_DM_WIDTH ( 4 ),
      .C_MIO_PRIMITIVE ( 54 ),
      .C_PACKAGE_NAME ( "clg484" ),
      .C_PS7_SI_REV ( "PRODUCTION" ),
      .C_M_AXI_GP0_ID_WIDTH ( 12 ),
      .C_M_AXI_GP0_ENABLE_STATIC_REMAP ( 0 ),
      .C_M_AXI_GP1_ID_WIDTH ( 12 ),
      .C_M_AXI_GP1_ENABLE_STATIC_REMAP ( 0 ),
      .C_S_AXI_GP0_ID_WIDTH ( 6 ),
      .C_S_AXI_GP1_ID_WIDTH ( 6 ),
      .C_S_AXI_ACP_ID_WIDTH ( 3 ),
      .C_S_AXI_HP0_ID_WIDTH ( 2 ),
      .C_S_AXI_HP0_DATA_WIDTH ( 64 ),
      .C_S_AXI_HP1_ID_WIDTH ( 6 ),
      .C_S_AXI_HP1_DATA_WIDTH ( 64 ),
      .C_S_AXI_HP2_ID_WIDTH ( 6 ),
      .C_S_AXI_HP2_DATA_WIDTH ( 64 ),
      .C_S_AXI_HP3_ID_WIDTH ( 6 ),
      .C_S_AXI_HP3_DATA_WIDTH ( 64 ),
      .C_M_AXI_GP0_THREAD_ID_WIDTH ( 12 ),
      .C_M_AXI_GP1_THREAD_ID_WIDTH ( 12 ),
      .C_NUM_F2P_INTR_INPUTS ( 1 ),
      .C_FCLK_CLK0_BUF ( "TRUE" ),
      .C_FCLK_CLK1_BUF ( "FALSE" ),
      .C_FCLK_CLK2_BUF ( "FALSE" ),
      .C_FCLK_CLK3_BUF ( "TRUE" )
    )
    processing_system7_0 (
      .CAN0_PHY_TX ( CAN0_PHY_TX ),
      .CAN0_PHY_RX ( CAN0_PHY_RX ),
      .CAN1_PHY_TX ( CAN1_PHY_TX ),
      .CAN1_PHY_RX ( CAN1_PHY_RX ),
      .ENET0_GMII_TX_EN ( ENET0_GMII_TX_EN ),
      .ENET0_GMII_TX_ER ( ENET0_GMII_TX_ER ),
      .ENET0_MDIO_MDC ( ENET0_MDIO_MDC ),
      .ENET0_MDIO_O ( ENET0_MDIO_O ),
      .ENET0_MDIO_T ( ENET0_MDIO_T ),
      .ENET0_PTP_DELAY_REQ_RX ( ENET0_PTP_DELAY_REQ_RX ),
      .ENET0_PTP_DELAY_REQ_TX ( ENET0_PTP_DELAY_REQ_TX ),
      .ENET0_PTP_PDELAY_REQ_RX ( ENET0_PTP_PDELAY_REQ_RX ),
      .ENET0_PTP_PDELAY_REQ_TX ( ENET0_PTP_PDELAY_REQ_TX ),
      .ENET0_PTP_PDELAY_RESP_RX ( ENET0_PTP_PDELAY_RESP_RX ),
      .ENET0_PTP_PDELAY_RESP_TX ( ENET0_PTP_PDELAY_RESP_TX ),
      .ENET0_PTP_SYNC_FRAME_RX ( ENET0_PTP_SYNC_FRAME_RX ),
      .ENET0_PTP_SYNC_FRAME_TX ( ENET0_PTP_SYNC_FRAME_TX ),
      .ENET0_SOF_RX ( ENET0_SOF_RX ),
      .ENET0_SOF_TX ( ENET0_SOF_TX ),
      .ENET0_GMII_TXD ( ENET0_GMII_TXD ),
      .ENET0_GMII_COL ( ENET0_GMII_COL ),
      .ENET0_GMII_CRS ( ENET0_GMII_CRS ),
      .ENET0_EXT_INTIN ( ENET0_EXT_INTIN ),
      .ENET0_GMII_RX_CLK ( ENET0_GMII_RX_CLK ),
      .ENET0_GMII_RX_DV ( ENET0_GMII_RX_DV ),
      .ENET0_GMII_RX_ER ( ENET0_GMII_RX_ER ),
      .ENET0_GMII_TX_CLK ( ENET0_GMII_TX_CLK ),
      .ENET0_MDIO_I ( ENET0_MDIO_I ),
      .ENET0_GMII_RXD ( ENET0_GMII_RXD ),
      .ENET1_GMII_TX_EN ( ENET1_GMII_TX_EN ),
      .ENET1_GMII_TX_ER ( ENET1_GMII_TX_ER ),
      .ENET1_MDIO_MDC ( ENET1_MDIO_MDC ),
      .ENET1_MDIO_O ( ENET1_MDIO_O ),
      .ENET1_MDIO_T ( ENET1_MDIO_T ),
      .ENET1_PTP_DELAY_REQ_RX ( ENET1_PTP_DELAY_REQ_RX ),
      .ENET1_PTP_DELAY_REQ_TX ( ENET1_PTP_DELAY_REQ_TX ),
      .ENET1_PTP_PDELAY_REQ_RX ( ENET1_PTP_PDELAY_REQ_RX ),
      .ENET1_PTP_PDELAY_REQ_TX ( ENET1_PTP_PDELAY_REQ_TX ),
      .ENET1_PTP_PDELAY_RESP_RX ( ENET1_PTP_PDELAY_RESP_RX ),
      .ENET1_PTP_PDELAY_RESP_TX ( ENET1_PTP_PDELAY_RESP_TX ),
      .ENET1_PTP_SYNC_FRAME_RX ( ENET1_PTP_SYNC_FRAME_RX ),
      .ENET1_PTP_SYNC_FRAME_TX ( ENET1_PTP_SYNC_FRAME_TX ),
      .ENET1_SOF_RX ( ENET1_SOF_RX ),
      .ENET1_SOF_TX ( ENET1_SOF_TX ),
      .ENET1_GMII_TXD ( ENET1_GMII_TXD ),
      .ENET1_GMII_COL ( ENET1_GMII_COL ),
      .ENET1_GMII_CRS ( ENET1_GMII_CRS ),
      .ENET1_EXT_INTIN ( ENET1_EXT_INTIN ),
      .ENET1_GMII_RX_CLK ( ENET1_GMII_RX_CLK ),
      .ENET1_GMII_RX_DV ( ENET1_GMII_RX_DV ),
      .ENET1_GMII_RX_ER ( ENET1_GMII_RX_ER ),
      .ENET1_GMII_TX_CLK ( ENET1_GMII_TX_CLK ),
      .ENET1_MDIO_I ( ENET1_MDIO_I ),
      .ENET1_GMII_RXD ( ENET1_GMII_RXD ),
      .GPIO_I ( GPIO_I ),
      .GPIO_O ( GPIO_O ),
      .GPIO_T ( GPIO_T ),
      .I2C0_SDA_I ( I2C0_SDA_I ),
      .I2C0_SDA_O ( I2C0_SDA_O ),
      .I2C0_SDA_T ( I2C0_SDA_T ),
      .I2C0_SCL_I ( I2C0_SCL_I ),
      .I2C0_SCL_O ( I2C0_SCL_O ),
      .I2C0_SCL_T ( I2C0_SCL_T ),
      .I2C1_SDA_I ( I2C1_SDA_I ),
      .I2C1_SDA_O ( I2C1_SDA_O ),
      .I2C1_SDA_T ( I2C1_SDA_T ),
      .I2C1_SCL_I ( I2C1_SCL_I ),
      .I2C1_SCL_O ( I2C1_SCL_O ),
      .I2C1_SCL_T ( I2C1_SCL_T ),
      .PJTAG_TCK ( PJTAG_TCK ),
      .PJTAG_TMS ( PJTAG_TMS ),
      .PJTAG_TD_I ( PJTAG_TD_I ),
      .PJTAG_TD_T ( PJTAG_TD_T ),
      .PJTAG_TD_O ( PJTAG_TD_O ),
      .SDIO0_CLK ( SDIO0_CLK ),
      .SDIO0_CLK_FB ( SDIO0_CLK_FB ),
      .SDIO0_CMD_O ( SDIO0_CMD_O ),
      .SDIO0_CMD_I ( SDIO0_CMD_I ),
      .SDIO0_CMD_T ( SDIO0_CMD_T ),
      .SDIO0_DATA_I ( SDIO0_DATA_I ),
      .SDIO0_DATA_O ( SDIO0_DATA_O ),
      .SDIO0_DATA_T ( SDIO0_DATA_T ),
      .SDIO0_LED ( SDIO0_LED ),
      .SDIO0_CDN ( SDIO0_CDN ),
      .SDIO0_WP ( SDIO0_WP ),
      .SDIO0_BUSPOW ( SDIO0_BUSPOW ),
      .SDIO0_BUSVOLT ( SDIO0_BUSVOLT ),
      .SDIO1_CLK ( SDIO1_CLK ),
      .SDIO1_CLK_FB ( SDIO1_CLK_FB ),
      .SDIO1_CMD_O ( SDIO1_CMD_O ),
      .SDIO1_CMD_I ( SDIO1_CMD_I ),
      .SDIO1_CMD_T ( SDIO1_CMD_T ),
      .SDIO1_DATA_I ( SDIO1_DATA_I ),
      .SDIO1_DATA_O ( SDIO1_DATA_O ),
      .SDIO1_DATA_T ( SDIO1_DATA_T ),
      .SDIO1_LED ( SDIO1_LED ),
      .SDIO1_CDN ( SDIO1_CDN ),
      .SDIO1_WP ( SDIO1_WP ),
      .SDIO1_BUSPOW ( SDIO1_BUSPOW ),
      .SDIO1_BUSVOLT ( SDIO1_BUSVOLT ),
      .SPI0_SCLK_I ( SPI0_SCLK_I ),
      .SPI0_SCLK_O ( SPI0_SCLK_O ),
      .SPI0_SCLK_T ( SPI0_SCLK_T ),
      .SPI0_MOSI_I ( SPI0_MOSI_I ),
      .SPI0_MOSI_O ( SPI0_MOSI_O ),
      .SPI0_MOSI_T ( SPI0_MOSI_T ),
      .SPI0_MISO_I ( SPI0_MISO_I ),
      .SPI0_MISO_O ( SPI0_MISO_O ),
      .SPI0_MISO_T ( SPI0_MISO_T ),
      .SPI0_SS_I ( SPI0_SS_I ),
      .SPI0_SS_O ( SPI0_SS_O ),
      .SPI0_SS1_O ( SPI0_SS1_O ),
      .SPI0_SS2_O ( SPI0_SS2_O ),
      .SPI0_SS_T ( SPI0_SS_T ),
      .SPI1_SCLK_I ( SPI1_SCLK_I ),
      .SPI1_SCLK_O ( SPI1_SCLK_O ),
      .SPI1_SCLK_T ( SPI1_SCLK_T ),
      .SPI1_MOSI_I ( SPI1_MOSI_I ),
      .SPI1_MOSI_O ( SPI1_MOSI_O ),
      .SPI1_MOSI_T ( SPI1_MOSI_T ),
      .SPI1_MISO_I ( SPI1_MISO_I ),
      .SPI1_MISO_O ( SPI1_MISO_O ),
      .SPI1_MISO_T ( SPI1_MISO_T ),
      .SPI1_SS_I ( SPI1_SS_I ),
      .SPI1_SS_O ( SPI1_SS_O ),
      .SPI1_SS1_O ( SPI1_SS1_O ),
      .SPI1_SS2_O ( SPI1_SS2_O ),
      .SPI1_SS_T ( SPI1_SS_T ),
      .UART0_DTRN ( UART0_DTRN ),
      .UART0_RTSN ( UART0_RTSN ),
      .UART0_TX ( UART0_TX ),
      .UART0_CTSN ( UART0_CTSN ),
      .UART0_DCDN ( UART0_DCDN ),
      .UART0_DSRN ( UART0_DSRN ),
      .UART0_RIN ( UART0_RIN ),
      .UART0_RX ( UART0_RX ),
      .UART1_DTRN ( UART1_DTRN ),
      .UART1_RTSN ( UART1_RTSN ),
      .UART1_TX ( UART1_TX ),
      .UART1_CTSN ( UART1_CTSN ),
      .UART1_DCDN ( UART1_DCDN ),
      .UART1_DSRN ( UART1_DSRN ),
      .UART1_RIN ( UART1_RIN ),
      .UART1_RX ( UART1_RX ),
      .TTC0_WAVE0_OUT ( TTC0_WAVE0_OUT ),
      .TTC0_WAVE1_OUT ( TTC0_WAVE1_OUT ),
      .TTC0_WAVE2_OUT ( TTC0_WAVE2_OUT ),
      .TTC0_CLK0_IN ( TTC0_CLK0_IN ),
      .TTC0_CLK1_IN ( TTC0_CLK1_IN ),
      .TTC0_CLK2_IN ( TTC0_CLK2_IN ),
      .TTC1_WAVE0_OUT ( TTC1_WAVE0_OUT ),
      .TTC1_WAVE1_OUT ( TTC1_WAVE1_OUT ),
      .TTC1_WAVE2_OUT ( TTC1_WAVE2_OUT ),
      .TTC1_CLK0_IN ( TTC1_CLK0_IN ),
      .TTC1_CLK1_IN ( TTC1_CLK1_IN ),
      .TTC1_CLK2_IN ( TTC1_CLK2_IN ),
      .WDT_CLK_IN ( WDT_CLK_IN ),
      .WDT_RST_OUT ( WDT_RST_OUT ),
      .TRACE_CLK ( TRACE_CLK ),
      .TRACE_CTL ( TRACE_CTL ),
      .TRACE_DATA ( TRACE_DATA ),
      .USB0_PORT_INDCTL ( USB0_PORT_INDCTL ),
      .USB1_PORT_INDCTL ( USB1_PORT_INDCTL ),
      .USB0_VBUS_PWRSELECT ( USB0_VBUS_PWRSELECT ),
      .USB1_VBUS_PWRSELECT ( USB1_VBUS_PWRSELECT ),
      .USB0_VBUS_PWRFAULT ( USB0_VBUS_PWRFAULT ),
      .USB1_VBUS_PWRFAULT ( USB1_VBUS_PWRFAULT ),
      .SRAM_INTIN ( SRAM_INTIN ),
      .M_AXI_GP0_ARESETN ( M_AXI_GP0_ARESETN ),
      .M_AXI_GP0_ARVALID ( M_AXI_GP0_ARVALID ),
      .M_AXI_GP0_AWVALID ( M_AXI_GP0_AWVALID ),
      .M_AXI_GP0_BREADY ( M_AXI_GP0_BREADY ),
      .M_AXI_GP0_RREADY ( M_AXI_GP0_RREADY ),
      .M_AXI_GP0_WLAST ( M_AXI_GP0_WLAST ),
      .M_AXI_GP0_WVALID ( M_AXI_GP0_WVALID ),
      .M_AXI_GP0_ARID ( M_AXI_GP0_ARID ),
      .M_AXI_GP0_AWID ( M_AXI_GP0_AWID ),
      .M_AXI_GP0_WID ( M_AXI_GP0_WID ),
      .M_AXI_GP0_ARBURST ( M_AXI_GP0_ARBURST ),
      .M_AXI_GP0_ARLOCK ( M_AXI_GP0_ARLOCK ),
      .M_AXI_GP0_ARSIZE ( M_AXI_GP0_ARSIZE ),
      .M_AXI_GP0_AWBURST ( M_AXI_GP0_AWBURST ),
      .M_AXI_GP0_AWLOCK ( M_AXI_GP0_AWLOCK ),
      .M_AXI_GP0_AWSIZE ( M_AXI_GP0_AWSIZE ),
      .M_AXI_GP0_ARPROT ( M_AXI_GP0_ARPROT ),
      .M_AXI_GP0_AWPROT ( M_AXI_GP0_AWPROT ),
      .M_AXI_GP0_ARADDR ( M_AXI_GP0_ARADDR ),
      .M_AXI_GP0_AWADDR ( M_AXI_GP0_AWADDR ),
      .M_AXI_GP0_WDATA ( M_AXI_GP0_WDATA ),
      .M_AXI_GP0_ARCACHE ( M_AXI_GP0_ARCACHE ),
      .M_AXI_GP0_ARLEN ( M_AXI_GP0_ARLEN ),
      .M_AXI_GP0_ARQOS ( M_AXI_GP0_ARQOS ),
      .M_AXI_GP0_AWCACHE ( M_AXI_GP0_AWCACHE ),
      .M_AXI_GP0_AWLEN ( M_AXI_GP0_AWLEN ),
      .M_AXI_GP0_AWQOS ( M_AXI_GP0_AWQOS ),
      .M_AXI_GP0_WSTRB ( M_AXI_GP0_WSTRB ),
      .M_AXI_GP0_ACLK ( M_AXI_GP0_ACLK ),
      .M_AXI_GP0_ARREADY ( M_AXI_GP0_ARREADY ),
      .M_AXI_GP0_AWREADY ( M_AXI_GP0_AWREADY ),
      .M_AXI_GP0_BVALID ( M_AXI_GP0_BVALID ),
      .M_AXI_GP0_RLAST ( M_AXI_GP0_RLAST ),
      .M_AXI_GP0_RVALID ( M_AXI_GP0_RVALID ),
      .M_AXI_GP0_WREADY ( M_AXI_GP0_WREADY ),
      .M_AXI_GP0_BID ( M_AXI_GP0_BID ),
      .M_AXI_GP0_RID ( M_AXI_GP0_RID ),
      .M_AXI_GP0_BRESP ( M_AXI_GP0_BRESP ),
      .M_AXI_GP0_RRESP ( M_AXI_GP0_RRESP ),
      .M_AXI_GP0_RDATA ( M_AXI_GP0_RDATA ),
      .M_AXI_GP1_ARESETN ( M_AXI_GP1_ARESETN ),
      .M_AXI_GP1_ARVALID ( M_AXI_GP1_ARVALID ),
      .M_AXI_GP1_AWVALID ( M_AXI_GP1_AWVALID ),
      .M_AXI_GP1_BREADY ( M_AXI_GP1_BREADY ),
      .M_AXI_GP1_RREADY ( M_AXI_GP1_RREADY ),
      .M_AXI_GP1_WLAST ( M_AXI_GP1_WLAST ),
      .M_AXI_GP1_WVALID ( M_AXI_GP1_WVALID ),
      .M_AXI_GP1_ARID ( M_AXI_GP1_ARID ),
      .M_AXI_GP1_AWID ( M_AXI_GP1_AWID ),
      .M_AXI_GP1_WID ( M_AXI_GP1_WID ),
      .M_AXI_GP1_ARBURST ( M_AXI_GP1_ARBURST ),
      .M_AXI_GP1_ARLOCK ( M_AXI_GP1_ARLOCK ),
      .M_AXI_GP1_ARSIZE ( M_AXI_GP1_ARSIZE ),
      .M_AXI_GP1_AWBURST ( M_AXI_GP1_AWBURST ),
      .M_AXI_GP1_AWLOCK ( M_AXI_GP1_AWLOCK ),
      .M_AXI_GP1_AWSIZE ( M_AXI_GP1_AWSIZE ),
      .M_AXI_GP1_ARPROT ( M_AXI_GP1_ARPROT ),
      .M_AXI_GP1_AWPROT ( M_AXI_GP1_AWPROT ),
      .M_AXI_GP1_ARADDR ( M_AXI_GP1_ARADDR ),
      .M_AXI_GP1_AWADDR ( M_AXI_GP1_AWADDR ),
      .M_AXI_GP1_WDATA ( M_AXI_GP1_WDATA ),
      .M_AXI_GP1_ARCACHE ( M_AXI_GP1_ARCACHE ),
      .M_AXI_GP1_ARLEN ( M_AXI_GP1_ARLEN ),
      .M_AXI_GP1_ARQOS ( M_AXI_GP1_ARQOS ),
      .M_AXI_GP1_AWCACHE ( M_AXI_GP1_AWCACHE ),
      .M_AXI_GP1_AWLEN ( M_AXI_GP1_AWLEN ),
      .M_AXI_GP1_AWQOS ( M_AXI_GP1_AWQOS ),
      .M_AXI_GP1_WSTRB ( M_AXI_GP1_WSTRB ),
      .M_AXI_GP1_ACLK ( M_AXI_GP1_ACLK ),
      .M_AXI_GP1_ARREADY ( M_AXI_GP1_ARREADY ),
      .M_AXI_GP1_AWREADY ( M_AXI_GP1_AWREADY ),
      .M_AXI_GP1_BVALID ( M_AXI_GP1_BVALID ),
      .M_AXI_GP1_RLAST ( M_AXI_GP1_RLAST ),
      .M_AXI_GP1_RVALID ( M_AXI_GP1_RVALID ),
      .M_AXI_GP1_WREADY ( M_AXI_GP1_WREADY ),
      .M_AXI_GP1_BID ( M_AXI_GP1_BID ),
      .M_AXI_GP1_RID ( M_AXI_GP1_RID ),
      .M_AXI_GP1_BRESP ( M_AXI_GP1_BRESP ),
      .M_AXI_GP1_RRESP ( M_AXI_GP1_RRESP ),
      .M_AXI_GP1_RDATA ( M_AXI_GP1_RDATA ),
      .S_AXI_GP0_ARESETN ( S_AXI_GP0_ARESETN ),
      .S_AXI_GP0_ARREADY ( S_AXI_GP0_ARREADY ),
      .S_AXI_GP0_AWREADY ( S_AXI_GP0_AWREADY ),
      .S_AXI_GP0_BVALID ( S_AXI_GP0_BVALID ),
      .S_AXI_GP0_RLAST ( S_AXI_GP0_RLAST ),
      .S_AXI_GP0_RVALID ( S_AXI_GP0_RVALID ),
      .S_AXI_GP0_WREADY ( S_AXI_GP0_WREADY ),
      .S_AXI_GP0_BRESP ( S_AXI_GP0_BRESP ),
      .S_AXI_GP0_RRESP ( S_AXI_GP0_RRESP ),
      .S_AXI_GP0_RDATA ( S_AXI_GP0_RDATA ),
      .S_AXI_GP0_BID ( S_AXI_GP0_BID ),
      .S_AXI_GP0_RID ( S_AXI_GP0_RID ),
      .S_AXI_GP0_ACLK ( S_AXI_GP0_ACLK ),
      .S_AXI_GP0_ARVALID ( S_AXI_GP0_ARVALID ),
      .S_AXI_GP0_AWVALID ( S_AXI_GP0_AWVALID ),
      .S_AXI_GP0_BREADY ( S_AXI_GP0_BREADY ),
      .S_AXI_GP0_RREADY ( S_AXI_GP0_RREADY ),
      .S_AXI_GP0_WLAST ( S_AXI_GP0_WLAST ),
      .S_AXI_GP0_WVALID ( S_AXI_GP0_WVALID ),
      .S_AXI_GP0_ARBURST ( S_AXI_GP0_ARBURST ),
      .S_AXI_GP0_ARLOCK ( S_AXI_GP0_ARLOCK ),
      .S_AXI_GP0_ARSIZE ( S_AXI_GP0_ARSIZE ),
      .S_AXI_GP0_AWBURST ( S_AXI_GP0_AWBURST ),
      .S_AXI_GP0_AWLOCK ( S_AXI_GP0_AWLOCK ),
      .S_AXI_GP0_AWSIZE ( S_AXI_GP0_AWSIZE ),
      .S_AXI_GP0_ARPROT ( S_AXI_GP0_ARPROT ),
      .S_AXI_GP0_AWPROT ( S_AXI_GP0_AWPROT ),
      .S_AXI_GP0_ARADDR ( S_AXI_GP0_ARADDR ),
      .S_AXI_GP0_AWADDR ( S_AXI_GP0_AWADDR ),
      .S_AXI_GP0_WDATA ( S_AXI_GP0_WDATA ),
      .S_AXI_GP0_ARCACHE ( S_AXI_GP0_ARCACHE ),
      .S_AXI_GP0_ARLEN ( S_AXI_GP0_ARLEN ),
      .S_AXI_GP0_ARQOS ( S_AXI_GP0_ARQOS ),
      .S_AXI_GP0_AWCACHE ( S_AXI_GP0_AWCACHE ),
      .S_AXI_GP0_AWLEN ( S_AXI_GP0_AWLEN ),
      .S_AXI_GP0_AWQOS ( S_AXI_GP0_AWQOS ),
      .S_AXI_GP0_WSTRB ( S_AXI_GP0_WSTRB ),
      .S_AXI_GP0_ARID ( S_AXI_GP0_ARID ),
      .S_AXI_GP0_AWID ( S_AXI_GP0_AWID ),
      .S_AXI_GP0_WID ( S_AXI_GP0_WID ),
      .S_AXI_GP1_ARESETN ( S_AXI_GP1_ARESETN ),
      .S_AXI_GP1_ARREADY ( S_AXI_GP1_ARREADY ),
      .S_AXI_GP1_AWREADY ( S_AXI_GP1_AWREADY ),
      .S_AXI_GP1_BVALID ( S_AXI_GP1_BVALID ),
      .S_AXI_GP1_RLAST ( S_AXI_GP1_RLAST ),
      .S_AXI_GP1_RVALID ( S_AXI_GP1_RVALID ),
      .S_AXI_GP1_WREADY ( S_AXI_GP1_WREADY ),
      .S_AXI_GP1_BRESP ( S_AXI_GP1_BRESP ),
      .S_AXI_GP1_RRESP ( S_AXI_GP1_RRESP ),
      .S_AXI_GP1_RDATA ( S_AXI_GP1_RDATA ),
      .S_AXI_GP1_BID ( S_AXI_GP1_BID ),
      .S_AXI_GP1_RID ( S_AXI_GP1_RID ),
      .S_AXI_GP1_ACLK ( S_AXI_GP1_ACLK ),
      .S_AXI_GP1_ARVALID ( S_AXI_GP1_ARVALID ),
      .S_AXI_GP1_AWVALID ( S_AXI_GP1_AWVALID ),
      .S_AXI_GP1_BREADY ( S_AXI_GP1_BREADY ),
      .S_AXI_GP1_RREADY ( S_AXI_GP1_RREADY ),
      .S_AXI_GP1_WLAST ( S_AXI_GP1_WLAST ),
      .S_AXI_GP1_WVALID ( S_AXI_GP1_WVALID ),
      .S_AXI_GP1_ARBURST ( S_AXI_GP1_ARBURST ),
      .S_AXI_GP1_ARLOCK ( S_AXI_GP1_ARLOCK ),
      .S_AXI_GP1_ARSIZE ( S_AXI_GP1_ARSIZE ),
      .S_AXI_GP1_AWBURST ( S_AXI_GP1_AWBURST ),
      .S_AXI_GP1_AWLOCK ( S_AXI_GP1_AWLOCK ),
      .S_AXI_GP1_AWSIZE ( S_AXI_GP1_AWSIZE ),
      .S_AXI_GP1_ARPROT ( S_AXI_GP1_ARPROT ),
      .S_AXI_GP1_AWPROT ( S_AXI_GP1_AWPROT ),
      .S_AXI_GP1_ARADDR ( S_AXI_GP1_ARADDR ),
      .S_AXI_GP1_AWADDR ( S_AXI_GP1_AWADDR ),
      .S_AXI_GP1_WDATA ( S_AXI_GP1_WDATA ),
      .S_AXI_GP1_ARCACHE ( S_AXI_GP1_ARCACHE ),
      .S_AXI_GP1_ARLEN ( S_AXI_GP1_ARLEN ),
      .S_AXI_GP1_ARQOS ( S_AXI_GP1_ARQOS ),
      .S_AXI_GP1_AWCACHE ( S_AXI_GP1_AWCACHE ),
      .S_AXI_GP1_AWLEN ( S_AXI_GP1_AWLEN ),
      .S_AXI_GP1_AWQOS ( S_AXI_GP1_AWQOS ),
      .S_AXI_GP1_WSTRB ( S_AXI_GP1_WSTRB ),
      .S_AXI_GP1_ARID ( S_AXI_GP1_ARID ),
      .S_AXI_GP1_AWID ( S_AXI_GP1_AWID ),
      .S_AXI_GP1_WID ( S_AXI_GP1_WID ),
      .S_AXI_ACP_ARESETN ( S_AXI_ACP_ARESETN ),
      .S_AXI_ACP_AWREADY ( S_AXI_ACP_AWREADY ),
      .S_AXI_ACP_ARREADY ( S_AXI_ACP_ARREADY ),
      .S_AXI_ACP_BVALID ( S_AXI_ACP_BVALID ),
      .S_AXI_ACP_RLAST ( S_AXI_ACP_RLAST ),
      .S_AXI_ACP_RVALID ( S_AXI_ACP_RVALID ),
      .S_AXI_ACP_WREADY ( S_AXI_ACP_WREADY ),
      .S_AXI_ACP_BRESP ( S_AXI_ACP_BRESP ),
      .S_AXI_ACP_RRESP ( S_AXI_ACP_RRESP ),
      .S_AXI_ACP_BID ( S_AXI_ACP_BID ),
      .S_AXI_ACP_RID ( S_AXI_ACP_RID ),
      .S_AXI_ACP_RDATA ( S_AXI_ACP_RDATA ),
      .S_AXI_ACP_ACLK ( S_AXI_ACP_ACLK ),
      .S_AXI_ACP_ARVALID ( S_AXI_ACP_ARVALID ),
      .S_AXI_ACP_AWVALID ( S_AXI_ACP_AWVALID ),
      .S_AXI_ACP_BREADY ( S_AXI_ACP_BREADY ),
      .S_AXI_ACP_RREADY ( S_AXI_ACP_RREADY ),
      .S_AXI_ACP_WLAST ( S_AXI_ACP_WLAST ),
      .S_AXI_ACP_WVALID ( S_AXI_ACP_WVALID ),
      .S_AXI_ACP_ARID ( S_AXI_ACP_ARID ),
      .S_AXI_ACP_ARPROT ( S_AXI_ACP_ARPROT ),
      .S_AXI_ACP_AWID ( S_AXI_ACP_AWID ),
      .S_AXI_ACP_AWPROT ( S_AXI_ACP_AWPROT ),
      .S_AXI_ACP_WID ( S_AXI_ACP_WID ),
      .S_AXI_ACP_ARADDR ( S_AXI_ACP_ARADDR ),
      .S_AXI_ACP_AWADDR ( S_AXI_ACP_AWADDR ),
      .S_AXI_ACP_ARCACHE ( S_AXI_ACP_ARCACHE ),
      .S_AXI_ACP_ARLEN ( S_AXI_ACP_ARLEN ),
      .S_AXI_ACP_ARQOS ( S_AXI_ACP_ARQOS ),
      .S_AXI_ACP_AWCACHE ( S_AXI_ACP_AWCACHE ),
      .S_AXI_ACP_AWLEN ( S_AXI_ACP_AWLEN ),
      .S_AXI_ACP_AWQOS ( S_AXI_ACP_AWQOS ),
      .S_AXI_ACP_ARBURST ( S_AXI_ACP_ARBURST ),
      .S_AXI_ACP_ARLOCK ( S_AXI_ACP_ARLOCK ),
      .S_AXI_ACP_ARSIZE ( S_AXI_ACP_ARSIZE ),
      .S_AXI_ACP_AWBURST ( S_AXI_ACP_AWBURST ),
      .S_AXI_ACP_AWLOCK ( S_AXI_ACP_AWLOCK ),
      .S_AXI_ACP_AWSIZE ( S_AXI_ACP_AWSIZE ),
      .S_AXI_ACP_ARUSER ( S_AXI_ACP_ARUSER ),
      .S_AXI_ACP_AWUSER ( S_AXI_ACP_AWUSER ),
      .S_AXI_ACP_WDATA ( S_AXI_ACP_WDATA ),
      .S_AXI_ACP_WSTRB ( S_AXI_ACP_WSTRB ),
      .S_AXI_HP0_ARESETN ( S_AXI_HP0_ARESETN ),
      .S_AXI_HP0_ARREADY ( S_AXI_HP0_ARREADY ),
      .S_AXI_HP0_AWREADY ( S_AXI_HP0_AWREADY ),
      .S_AXI_HP0_BVALID ( S_AXI_HP0_BVALID ),
      .S_AXI_HP0_RLAST ( S_AXI_HP0_RLAST ),
      .S_AXI_HP0_RVALID ( S_AXI_HP0_RVALID ),
      .S_AXI_HP0_WREADY ( S_AXI_HP0_WREADY ),
      .S_AXI_HP0_BRESP ( S_AXI_HP0_BRESP ),
      .S_AXI_HP0_RRESP ( S_AXI_HP0_RRESP ),
      .S_AXI_HP0_BID ( S_AXI_HP0_BID ),
      .S_AXI_HP0_RID ( S_AXI_HP0_RID ),
      .S_AXI_HP0_RDATA ( S_AXI_HP0_RDATA ),
      .S_AXI_HP0_RCOUNT ( S_AXI_HP0_RCOUNT ),
      .S_AXI_HP0_WCOUNT ( S_AXI_HP0_WCOUNT ),
      .S_AXI_HP0_RACOUNT ( S_AXI_HP0_RACOUNT ),
      .S_AXI_HP0_WACOUNT ( S_AXI_HP0_WACOUNT ),
      .S_AXI_HP0_ACLK ( S_AXI_HP0_ACLK ),
      .S_AXI_HP0_ARVALID ( S_AXI_HP0_ARVALID ),
      .S_AXI_HP0_AWVALID ( S_AXI_HP0_AWVALID ),
      .S_AXI_HP0_BREADY ( S_AXI_HP0_BREADY ),
      .S_AXI_HP0_RDISSUECAP1_EN ( S_AXI_HP0_RDISSUECAP1_EN ),
      .S_AXI_HP0_RREADY ( S_AXI_HP0_RREADY ),
      .S_AXI_HP0_WLAST ( S_AXI_HP0_WLAST ),
      .S_AXI_HP0_WRISSUECAP1_EN ( S_AXI_HP0_WRISSUECAP1_EN ),
      .S_AXI_HP0_WVALID ( S_AXI_HP0_WVALID ),
      .S_AXI_HP0_ARBURST ( S_AXI_HP0_ARBURST ),
      .S_AXI_HP0_ARLOCK ( S_AXI_HP0_ARLOCK ),
      .S_AXI_HP0_ARSIZE ( S_AXI_HP0_ARSIZE ),
      .S_AXI_HP0_AWBURST ( S_AXI_HP0_AWBURST ),
      .S_AXI_HP0_AWLOCK ( S_AXI_HP0_AWLOCK ),
      .S_AXI_HP0_AWSIZE ( S_AXI_HP0_AWSIZE ),
      .S_AXI_HP0_ARPROT ( S_AXI_HP0_ARPROT ),
      .S_AXI_HP0_AWPROT ( S_AXI_HP0_AWPROT ),
      .S_AXI_HP0_ARADDR ( S_AXI_HP0_ARADDR ),
      .S_AXI_HP0_AWADDR ( S_AXI_HP0_AWADDR ),
      .S_AXI_HP0_ARCACHE ( S_AXI_HP0_ARCACHE ),
      .S_AXI_HP0_ARLEN ( S_AXI_HP0_ARLEN ),
      .S_AXI_HP0_ARQOS ( S_AXI_HP0_ARQOS ),
      .S_AXI_HP0_AWCACHE ( S_AXI_HP0_AWCACHE ),
      .S_AXI_HP0_AWLEN ( S_AXI_HP0_AWLEN ),
      .S_AXI_HP0_AWQOS ( S_AXI_HP0_AWQOS ),
      .S_AXI_HP0_ARID ( S_AXI_HP0_ARID ),
      .S_AXI_HP0_AWID ( S_AXI_HP0_AWID ),
      .S_AXI_HP0_WID ( S_AXI_HP0_WID ),
      .S_AXI_HP0_WDATA ( S_AXI_HP0_WDATA ),
      .S_AXI_HP0_WSTRB ( S_AXI_HP0_WSTRB ),
      .S_AXI_HP1_ARESETN ( S_AXI_HP1_ARESETN ),
      .S_AXI_HP1_ARREADY ( S_AXI_HP1_ARREADY ),
      .S_AXI_HP1_AWREADY ( S_AXI_HP1_AWREADY ),
      .S_AXI_HP1_BVALID ( S_AXI_HP1_BVALID ),
      .S_AXI_HP1_RLAST ( S_AXI_HP1_RLAST ),
      .S_AXI_HP1_RVALID ( S_AXI_HP1_RVALID ),
      .S_AXI_HP1_WREADY ( S_AXI_HP1_WREADY ),
      .S_AXI_HP1_BRESP ( S_AXI_HP1_BRESP ),
      .S_AXI_HP1_RRESP ( S_AXI_HP1_RRESP ),
      .S_AXI_HP1_BID ( S_AXI_HP1_BID ),
      .S_AXI_HP1_RID ( S_AXI_HP1_RID ),
      .S_AXI_HP1_RDATA ( S_AXI_HP1_RDATA ),
      .S_AXI_HP1_RCOUNT ( S_AXI_HP1_RCOUNT ),
      .S_AXI_HP1_WCOUNT ( S_AXI_HP1_WCOUNT ),
      .S_AXI_HP1_RACOUNT ( S_AXI_HP1_RACOUNT ),
      .S_AXI_HP1_WACOUNT ( S_AXI_HP1_WACOUNT ),
      .S_AXI_HP1_ACLK ( S_AXI_HP1_ACLK ),
      .S_AXI_HP1_ARVALID ( S_AXI_HP1_ARVALID ),
      .S_AXI_HP1_AWVALID ( S_AXI_HP1_AWVALID ),
      .S_AXI_HP1_BREADY ( S_AXI_HP1_BREADY ),
      .S_AXI_HP1_RDISSUECAP1_EN ( S_AXI_HP1_RDISSUECAP1_EN ),
      .S_AXI_HP1_RREADY ( S_AXI_HP1_RREADY ),
      .S_AXI_HP1_WLAST ( S_AXI_HP1_WLAST ),
      .S_AXI_HP1_WRISSUECAP1_EN ( S_AXI_HP1_WRISSUECAP1_EN ),
      .S_AXI_HP1_WVALID ( S_AXI_HP1_WVALID ),
      .S_AXI_HP1_ARBURST ( S_AXI_HP1_ARBURST ),
      .S_AXI_HP1_ARLOCK ( S_AXI_HP1_ARLOCK ),
      .S_AXI_HP1_ARSIZE ( S_AXI_HP1_ARSIZE ),
      .S_AXI_HP1_AWBURST ( S_AXI_HP1_AWBURST ),
      .S_AXI_HP1_AWLOCK ( S_AXI_HP1_AWLOCK ),
      .S_AXI_HP1_AWSIZE ( S_AXI_HP1_AWSIZE ),
      .S_AXI_HP1_ARPROT ( S_AXI_HP1_ARPROT ),
      .S_AXI_HP1_AWPROT ( S_AXI_HP1_AWPROT ),
      .S_AXI_HP1_ARADDR ( S_AXI_HP1_ARADDR ),
      .S_AXI_HP1_AWADDR ( S_AXI_HP1_AWADDR ),
      .S_AXI_HP1_ARCACHE ( S_AXI_HP1_ARCACHE ),
      .S_AXI_HP1_ARLEN ( S_AXI_HP1_ARLEN ),
      .S_AXI_HP1_ARQOS ( S_AXI_HP1_ARQOS ),
      .S_AXI_HP1_AWCACHE ( S_AXI_HP1_AWCACHE ),
      .S_AXI_HP1_AWLEN ( S_AXI_HP1_AWLEN ),
      .S_AXI_HP1_AWQOS ( S_AXI_HP1_AWQOS ),
      .S_AXI_HP1_ARID ( S_AXI_HP1_ARID ),
      .S_AXI_HP1_AWID ( S_AXI_HP1_AWID ),
      .S_AXI_HP1_WID ( S_AXI_HP1_WID ),
      .S_AXI_HP1_WDATA ( S_AXI_HP1_WDATA ),
      .S_AXI_HP1_WSTRB ( S_AXI_HP1_WSTRB ),
      .S_AXI_HP2_ARESETN ( S_AXI_HP2_ARESETN ),
      .S_AXI_HP2_ARREADY ( S_AXI_HP2_ARREADY ),
      .S_AXI_HP2_AWREADY ( S_AXI_HP2_AWREADY ),
      .S_AXI_HP2_BVALID ( S_AXI_HP2_BVALID ),
      .S_AXI_HP2_RLAST ( S_AXI_HP2_RLAST ),
      .S_AXI_HP2_RVALID ( S_AXI_HP2_RVALID ),
      .S_AXI_HP2_WREADY ( S_AXI_HP2_WREADY ),
      .S_AXI_HP2_BRESP ( S_AXI_HP2_BRESP ),
      .S_AXI_HP2_RRESP ( S_AXI_HP2_RRESP ),
      .S_AXI_HP2_BID ( S_AXI_HP2_BID ),
      .S_AXI_HP2_RID ( S_AXI_HP2_RID ),
      .S_AXI_HP2_RDATA ( S_AXI_HP2_RDATA ),
      .S_AXI_HP2_RCOUNT ( S_AXI_HP2_RCOUNT ),
      .S_AXI_HP2_WCOUNT ( S_AXI_HP2_WCOUNT ),
      .S_AXI_HP2_RACOUNT ( S_AXI_HP2_RACOUNT ),
      .S_AXI_HP2_WACOUNT ( S_AXI_HP2_WACOUNT ),
      .S_AXI_HP2_ACLK ( S_AXI_HP2_ACLK ),
      .S_AXI_HP2_ARVALID ( S_AXI_HP2_ARVALID ),
      .S_AXI_HP2_AWVALID ( S_AXI_HP2_AWVALID ),
      .S_AXI_HP2_BREADY ( S_AXI_HP2_BREADY ),
      .S_AXI_HP2_RDISSUECAP1_EN ( S_AXI_HP2_RDISSUECAP1_EN ),
      .S_AXI_HP2_RREADY ( S_AXI_HP2_RREADY ),
      .S_AXI_HP2_WLAST ( S_AXI_HP2_WLAST ),
      .S_AXI_HP2_WRISSUECAP1_EN ( S_AXI_HP2_WRISSUECAP1_EN ),
      .S_AXI_HP2_WVALID ( S_AXI_HP2_WVALID ),
      .S_AXI_HP2_ARBURST ( S_AXI_HP2_ARBURST ),
      .S_AXI_HP2_ARLOCK ( S_AXI_HP2_ARLOCK ),
      .S_AXI_HP2_ARSIZE ( S_AXI_HP2_ARSIZE ),
      .S_AXI_HP2_AWBURST ( S_AXI_HP2_AWBURST ),
      .S_AXI_HP2_AWLOCK ( S_AXI_HP2_AWLOCK ),
      .S_AXI_HP2_AWSIZE ( S_AXI_HP2_AWSIZE ),
      .S_AXI_HP2_ARPROT ( S_AXI_HP2_ARPROT ),
      .S_AXI_HP2_AWPROT ( S_AXI_HP2_AWPROT ),
      .S_AXI_HP2_ARADDR ( S_AXI_HP2_ARADDR ),
      .S_AXI_HP2_AWADDR ( S_AXI_HP2_AWADDR ),
      .S_AXI_HP2_ARCACHE ( S_AXI_HP2_ARCACHE ),
      .S_AXI_HP2_ARLEN ( S_AXI_HP2_ARLEN ),
      .S_AXI_HP2_ARQOS ( S_AXI_HP2_ARQOS ),
      .S_AXI_HP2_AWCACHE ( S_AXI_HP2_AWCACHE ),
      .S_AXI_HP2_AWLEN ( S_AXI_HP2_AWLEN ),
      .S_AXI_HP2_AWQOS ( S_AXI_HP2_AWQOS ),
      .S_AXI_HP2_ARID ( S_AXI_HP2_ARID ),
      .S_AXI_HP2_AWID ( S_AXI_HP2_AWID ),
      .S_AXI_HP2_WID ( S_AXI_HP2_WID ),
      .S_AXI_HP2_WDATA ( S_AXI_HP2_WDATA ),
      .S_AXI_HP2_WSTRB ( S_AXI_HP2_WSTRB ),
      .S_AXI_HP3_ARESETN ( S_AXI_HP3_ARESETN ),
      .S_AXI_HP3_ARREADY ( S_AXI_HP3_ARREADY ),
      .S_AXI_HP3_AWREADY ( S_AXI_HP3_AWREADY ),
      .S_AXI_HP3_BVALID ( S_AXI_HP3_BVALID ),
      .S_AXI_HP3_RLAST ( S_AXI_HP3_RLAST ),
      .S_AXI_HP3_RVALID ( S_AXI_HP3_RVALID ),
      .S_AXI_HP3_WREADY ( S_AXI_HP3_WREADY ),
      .S_AXI_HP3_BRESP ( S_AXI_HP3_BRESP ),
      .S_AXI_HP3_RRESP ( S_AXI_HP3_RRESP ),
      .S_AXI_HP3_BID ( S_AXI_HP3_BID ),
      .S_AXI_HP3_RID ( S_AXI_HP3_RID ),
      .S_AXI_HP3_RDATA ( S_AXI_HP3_RDATA ),
      .S_AXI_HP3_RCOUNT ( S_AXI_HP3_RCOUNT ),
      .S_AXI_HP3_WCOUNT ( S_AXI_HP3_WCOUNT ),
      .S_AXI_HP3_RACOUNT ( S_AXI_HP3_RACOUNT ),
      .S_AXI_HP3_WACOUNT ( S_AXI_HP3_WACOUNT ),
      .S_AXI_HP3_ACLK ( S_AXI_HP3_ACLK ),
      .S_AXI_HP3_ARVALID ( S_AXI_HP3_ARVALID ),
      .S_AXI_HP3_AWVALID ( S_AXI_HP3_AWVALID ),
      .S_AXI_HP3_BREADY ( S_AXI_HP3_BREADY ),
      .S_AXI_HP3_RDISSUECAP1_EN ( S_AXI_HP3_RDISSUECAP1_EN ),
      .S_AXI_HP3_RREADY ( S_AXI_HP3_RREADY ),
      .S_AXI_HP3_WLAST ( S_AXI_HP3_WLAST ),
      .S_AXI_HP3_WRISSUECAP1_EN ( S_AXI_HP3_WRISSUECAP1_EN ),
      .S_AXI_HP3_WVALID ( S_AXI_HP3_WVALID ),
      .S_AXI_HP3_ARBURST ( S_AXI_HP3_ARBURST ),
      .S_AXI_HP3_ARLOCK ( S_AXI_HP3_ARLOCK ),
      .S_AXI_HP3_ARSIZE ( S_AXI_HP3_ARSIZE ),
      .S_AXI_HP3_AWBURST ( S_AXI_HP3_AWBURST ),
      .S_AXI_HP3_AWLOCK ( S_AXI_HP3_AWLOCK ),
      .S_AXI_HP3_AWSIZE ( S_AXI_HP3_AWSIZE ),
      .S_AXI_HP3_ARPROT ( S_AXI_HP3_ARPROT ),
      .S_AXI_HP3_AWPROT ( S_AXI_HP3_AWPROT ),
      .S_AXI_HP3_ARADDR ( S_AXI_HP3_ARADDR ),
      .S_AXI_HP3_AWADDR ( S_AXI_HP3_AWADDR ),
      .S_AXI_HP3_ARCACHE ( S_AXI_HP3_ARCACHE ),
      .S_AXI_HP3_ARLEN ( S_AXI_HP3_ARLEN ),
      .S_AXI_HP3_ARQOS ( S_AXI_HP3_ARQOS ),
      .S_AXI_HP3_AWCACHE ( S_AXI_HP3_AWCACHE ),
      .S_AXI_HP3_AWLEN ( S_AXI_HP3_AWLEN ),
      .S_AXI_HP3_AWQOS ( S_AXI_HP3_AWQOS ),
      .S_AXI_HP3_ARID ( S_AXI_HP3_ARID ),
      .S_AXI_HP3_AWID ( S_AXI_HP3_AWID ),
      .S_AXI_HP3_WID ( S_AXI_HP3_WID ),
      .S_AXI_HP3_WDATA ( S_AXI_HP3_WDATA ),
      .S_AXI_HP3_WSTRB ( S_AXI_HP3_WSTRB ),
      .DMA0_DATYPE ( DMA0_DATYPE ),
      .DMA0_DAVALID ( DMA0_DAVALID ),
      .DMA0_DRREADY ( DMA0_DRREADY ),
      .DMA0_RSTN ( DMA0_RSTN ),
      .DMA0_ACLK ( DMA0_ACLK ),
      .DMA0_DAREADY ( DMA0_DAREADY ),
      .DMA0_DRLAST ( DMA0_DRLAST ),
      .DMA0_DRVALID ( DMA0_DRVALID ),
      .DMA0_DRTYPE ( DMA0_DRTYPE ),
      .DMA1_DATYPE ( DMA1_DATYPE ),
      .DMA1_DAVALID ( DMA1_DAVALID ),
      .DMA1_DRREADY ( DMA1_DRREADY ),
      .DMA1_RSTN ( DMA1_RSTN ),
      .DMA1_ACLK ( DMA1_ACLK ),
      .DMA1_DAREADY ( DMA1_DAREADY ),
      .DMA1_DRLAST ( DMA1_DRLAST ),
      .DMA1_DRVALID ( DMA1_DRVALID ),
      .DMA1_DRTYPE ( DMA1_DRTYPE ),
      .DMA2_DATYPE ( DMA2_DATYPE ),
      .DMA2_DAVALID ( DMA2_DAVALID ),
      .DMA2_DRREADY ( DMA2_DRREADY ),
      .DMA2_RSTN ( DMA2_RSTN ),
      .DMA2_ACLK ( DMA2_ACLK ),
      .DMA2_DAREADY ( DMA2_DAREADY ),
      .DMA2_DRLAST ( DMA2_DRLAST ),
      .DMA2_DRVALID ( DMA2_DRVALID ),
      .DMA3_DRVALID ( DMA3_DRVALID ),
      .DMA3_DATYPE ( DMA3_DATYPE ),
      .DMA3_DAVALID ( DMA3_DAVALID ),
      .DMA3_DRREADY ( DMA3_DRREADY ),
      .DMA3_RSTN ( DMA3_RSTN ),
      .DMA3_ACLK ( DMA3_ACLK ),
      .DMA3_DAREADY ( DMA3_DAREADY ),
      .DMA3_DRLAST ( DMA3_DRLAST ),
      .DMA2_DRTYPE ( DMA2_DRTYPE ),
      .DMA3_DRTYPE ( DMA3_DRTYPE ),
      .FTMD_TRACEIN_DATA ( FTMD_TRACEIN_DATA ),
      .FTMD_TRACEIN_VALID ( FTMD_TRACEIN_VALID ),
      .FTMD_TRACEIN_CLK ( FTMD_TRACEIN_CLK ),
      .FTMD_TRACEIN_ATID ( FTMD_TRACEIN_ATID ),
      .FTMT_F2P_TRIG ( FTMT_F2P_TRIG ),
      .FTMT_F2P_TRIGACK ( FTMT_F2P_TRIGACK ),
      .FTMT_F2P_DEBUG ( FTMT_F2P_DEBUG ),
      .FTMT_P2F_TRIGACK ( FTMT_P2F_TRIGACK ),
      .FTMT_P2F_TRIG ( FTMT_P2F_TRIG ),
      .FTMT_P2F_DEBUG ( FTMT_P2F_DEBUG ),
      .FCLK_CLK3 ( FCLK_CLK3 ),
      .FCLK_CLK2 ( FCLK_CLK2 ),
      .FCLK_CLK1 ( FCLK_CLK1 ),
      .FCLK_CLK0 ( FCLK_CLK0 ),
      .FCLK_CLKTRIG3_N ( FCLK_CLKTRIG3_N ),
      .FCLK_CLKTRIG2_N ( FCLK_CLKTRIG2_N ),
      .FCLK_CLKTRIG1_N ( FCLK_CLKTRIG1_N ),
      .FCLK_CLKTRIG0_N ( FCLK_CLKTRIG0_N ),
      .FCLK_RESET3_N ( FCLK_RESET3_N ),
      .FCLK_RESET2_N ( FCLK_RESET2_N ),
      .FCLK_RESET1_N ( FCLK_RESET1_N ),
      .FCLK_RESET0_N ( FCLK_RESET0_N ),
      .FPGA_IDLE_N ( FPGA_IDLE_N ),
      .DDR_ARB ( DDR_ARB ),
      .IRQ_F2P ( IRQ_F2P ),
      .Core0_nFIQ ( Core0_nFIQ ),
      .Core0_nIRQ ( Core0_nIRQ ),
      .Core1_nFIQ ( Core1_nFIQ ),
      .Core1_nIRQ ( Core1_nIRQ ),
      .EVENT_EVENTO ( EVENT_EVENTO ),
      .EVENT_STANDBYWFE ( EVENT_STANDBYWFE ),
      .EVENT_STANDBYWFI ( EVENT_STANDBYWFI ),
      .EVENT_EVENTI ( EVENT_EVENTI ),
      .MIO ( MIO ),
      .DDR_Clk ( DDR_Clk ),
      .DDR_Clk_n ( DDR_Clk_n ),
      .DDR_CKE ( DDR_CKE ),
      .DDR_CS_n ( DDR_CS_n ),
      .DDR_RAS_n ( DDR_RAS_n ),
      .DDR_CAS_n ( DDR_CAS_n ),
      .DDR_WEB ( DDR_WEB ),
      .DDR_BankAddr ( DDR_BankAddr ),
      .DDR_Addr ( DDR_Addr ),
      .DDR_ODT ( DDR_ODT ),
      .DDR_DRSTB ( DDR_DRSTB ),
      .DDR_DQ ( DDR_DQ ),
      .DDR_DM ( DDR_DM ),
      .DDR_DQS ( DDR_DQS ),
      .DDR_DQS_n ( DDR_DQS_n ),
      .DDR_VRN ( DDR_VRN ),
      .DDR_VRP ( DDR_VRP ),
      .PS_SRSTB ( PS_SRSTB ),
      .PS_CLK ( PS_CLK ),
      .PS_PORB ( PS_PORB ),
      .IRQ_P2F_DMAC_ABORT ( IRQ_P2F_DMAC_ABORT ),
      .IRQ_P2F_DMAC0 ( IRQ_P2F_DMAC0 ),
      .IRQ_P2F_DMAC1 ( IRQ_P2F_DMAC1 ),
      .IRQ_P2F_DMAC2 ( IRQ_P2F_DMAC2 ),
      .IRQ_P2F_DMAC3 ( IRQ_P2F_DMAC3 ),
      .IRQ_P2F_DMAC4 ( IRQ_P2F_DMAC4 ),
      .IRQ_P2F_DMAC5 ( IRQ_P2F_DMAC5 ),
      .IRQ_P2F_DMAC6 ( IRQ_P2F_DMAC6 ),
      .IRQ_P2F_DMAC7 ( IRQ_P2F_DMAC7 ),
      .IRQ_P2F_SMC ( IRQ_P2F_SMC ),
      .IRQ_P2F_QSPI ( IRQ_P2F_QSPI ),
      .IRQ_P2F_CTI ( IRQ_P2F_CTI ),
      .IRQ_P2F_GPIO ( IRQ_P2F_GPIO ),
      .IRQ_P2F_USB0 ( IRQ_P2F_USB0 ),
      .IRQ_P2F_ENET0 ( IRQ_P2F_ENET0 ),
      .IRQ_P2F_ENET_WAKE0 ( IRQ_P2F_ENET_WAKE0 ),
      .IRQ_P2F_SDIO0 ( IRQ_P2F_SDIO0 ),
      .IRQ_P2F_I2C0 ( IRQ_P2F_I2C0 ),
      .IRQ_P2F_SPI0 ( IRQ_P2F_SPI0 ),
      .IRQ_P2F_UART0 ( IRQ_P2F_UART0 ),
      .IRQ_P2F_CAN0 ( IRQ_P2F_CAN0 ),
      .IRQ_P2F_USB1 ( IRQ_P2F_USB1 ),
      .IRQ_P2F_ENET1 ( IRQ_P2F_ENET1 ),
      .IRQ_P2F_ENET_WAKE1 ( IRQ_P2F_ENET_WAKE1 ),
      .IRQ_P2F_SDIO1 ( IRQ_P2F_SDIO1 ),
      .IRQ_P2F_I2C1 ( IRQ_P2F_I2C1 ),
      .IRQ_P2F_SPI1 ( IRQ_P2F_SPI1 ),
      .IRQ_P2F_UART1 ( IRQ_P2F_UART1 ),
      .IRQ_P2F_CAN1 ( IRQ_P2F_CAN1 )
    );

endmodule

