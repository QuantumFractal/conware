XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��w�=��D�&n/N�G!���Ajx��������K�!��l���%�-X�9M�6|;7��+X	9��i���E�?኉Q-�_m��y�@<J�������(E���n�/�:1T��_K]�l+zB+�N�)H���\,
��p��Ȋ�L�jӚOƮ���%C�]���w���J�?�Y3홤s�dL$�DŨ.�5�H�4/z���2L�+F,l�(�ϕu MK��I^�L�ґ�7��4K�~R��0�Ӫ؊N�����>�q�i�=Q4n��]�`O�tR�����<��lR	�!m��َKE�E@?�(��u$�:��Kh��60�
�֩,�CTY����\z�P�y�)�U��S�H�+1�ha�K�e��&$��%3h4IB*�lh3��x%�VT�s9��V�&���pF��3݆�b�K\�T���:ΎIt%p]���m���EŐ#���;{:�E��.�2]C��(���f�sٟ�u���T8�����&�K5��1�g�G%im�k��'��UH�B{p�JkǺrb�͒��{����ڽ��6*�8�ǡ9�a���A�\��l��M�9톡��Vo�"�b����B��HK���>�f�БY_2�$=/d�H(%��_��,������J�j�]��+�I���Y��߇��>,��[��O�~$��	]~�9%ob�k�����s�D\��q2X���H
��}�S!���B�Ӑ���ߜ������Q�S��(��;|�h���U��&�XlxVHYEB    3fdc    1160
x$�'M����j���
^�
��"7R*g��\
��]ߚW?�h���)�DB�T�0�YQe4�:1:�TL�<�:Z�Ι�#]��!lqli�_rs��r���M����:��,z��C�� U��ɩd���c��6EEwA��aݝxw��W�_�[[m�o���� �^%3��&��.�[j����+��9��@D�@�:������s���;���@��.��wv�b�3��͵��z�(wS����8��`�
m�/_�b��~"�Ww p�/���KDz![��C�	M�L�dG'��yP�	eD�׷b��N����3�XME��m�}G:�z�&�]�s�&9E���X�=j��aE�d�?[ò�2�￻I��B[q��N=_�쨞e0�����9�?�$�QB5禟���/ ��~� �3/�Y�6ڄ0�;���Wٚ�C:.l���ߋ����y�c�G�ʼ��~�	����+�X�Xm{�,���
a�f�J�5$�d�w�l�)���,`@K(=R���n�T�:�@��(�,��1��!(&篁�K���j*�&q���)���/R@<�$���Y)�\ �#���H�g��p�Z��@J\�-p�z�Y�Nދo��)�T���d���x<+!��[��R
X��
E�&���������*�!��Z�_�2PL��JXo�2���h��Ic����d��W���
2k�����r�;�<�E|���������#���&�Z���[��&G���sv�8Vk�?S�|Y;>�������p���~�e��<��;� ncl�f?ls�Xb���B�F?ف}
��j�L����<����T������ |�Շ�r��M����I~���+�j��.>s^�)u���zN�����y0;0*�����8�x��}CsK��hyL{]֐hAa<PSg���bJ�2;��A�r�'ڟ�/�����F����CRô�SK�4Mg���Ă����v2�1yTn�6�6]n�yhl�8�� _��
����v����T	o C�_k�D\c�&�M_�����B"p��܁^�]5S�~�H�ʁt�~�!����'F:ϛ�����N�V��c(�h	N���˟����7�~���.CȤ���"�y�/Z�o�-'{�m�H�E[���j�G�2��q ��&MS�M���H��6?w騉� p"#��aݩ�m'D@7\s�|���������M�<�Y3�1eyp�4�e)�%ם��@�ڭ������-X`��JM����ҫ>u��q�]l�軒[7������+�V����B>a��I#E&R�ôₔݽR8׿e�^*�I���"u�N,��%���n&T?��l�a��ގ���)�IQ��e��UR��y��L����Z�f�N�;�ܲ�+Y S�d��ƨ�n��^��l�;�3�{.�`�:�ˍ}��9�T�%�������ԋ��])�X�����sې�@������=��]/�V���ҎNJ�%hR�Ia��~���
�S\y��84�=�PT��à�Y<��@����x�o(���Ǆ�f�ڠXP#Tn��Nb�sV�"a�`,*���g�>�d�|��-$��پ��|�����(@i;6��
�Ͼ| X�"�k�R��y ]� ������y�un�}����2���ےG���Q��ѐb��]�i�U�\/���<� ��-}���b�P���X�pg���+��\�wnh�v��� �{��r��	�$���G@�R��u�(����8����<������~]�Zz�NV�L����Gz�:��vlп4��^�?v����H�B�{T>�N6@��y �PZ�E��G7��0�9o�V('|�O:��L��~9�em�]-��T]-�%b�$~�j���tny+k<���+�{�>^*�d��Zyz��!�����s &�����C��d���>NY7Um�Ok��� �#��z�e�=��ݝ�}���=���ر~O2�w�������d:Db�]�н�\�sۋ���9݉�gʯ������^E�\x���u7I�+f#�����#�xڔ/E&u[ޡ�˂�擘�t�>�(�	F줮G�GH�O��Wnx��m�i�-	*@{��`5	c��e�mWs���v��D�-ˮ��
�AT�N	����P�v�ʬ�qe^ϰ���F���L��S�ݚ���&W3U���BU?���JdV�ܱ��y*Qz[Z��J��P��;tٳ�E�Y�����w3����{�o��Z����ǿ������E��o�q���$3D���j��Z=�*�ke}4�	�	*�BI���
B5���wῬR�a��>�2��Wo��um,���؍(�3z&Ȧb@��h#>Y���Xq	�p����Dۏ��Kp�*ΓJ����	򿖟��u��CFD^
�4��/4����G�w���k�ѡ�R9_\���0�N�d�P��Z7��7<d�$TI�:�&gμ@�TF딼�8(s����~����FdJ���,�fy�(��?ˊ�������w�W����j8�G;zX
�-�0zL6�9O��[I�UբDC�L7��j��K�ևҭ�Hm�������t�O}$�����ϛk��8�Pr솉8P�m�`�3"�N0�:�R�+|[�l�<�t4�7���݌�+���_k�a=g=��|�/�o̬��%�n�-��G�����/���9}�G�YDd�G��0�8^U�6�2y�$>L��Ĕ���@˳?�!|��ul�C��Q�p�K��,ղ��P��(�I�mf�o��-�� O�o�#9�*�d������됗�����
)�A�<���L�� �*����A�L�������f��҂d�U�j](��ϻ��T�z��8�#�{���[MJ�,4�$	��cd�Mml��T�v��m~<~7�M% �~O��y�9c@�=�T�`�����mY��v�Nk��y�~3k���&����(�,����A��g��zq�`��tG�������-�[)Δ3�� sGؐ��if8r ��$�}P�_����& ���pB� ˊrκ�G&��Y[�����=�(��p���fb_y�fϗ�o���F���R��uP�Lz-��/�L��:&��R�е�,�^������<��=V)�A�ɹ�`ջ�Y��b��{�y$/�!!�9v�`�g���RHZ�1�;:x�&�P�]S��/�[Q���T��(~`�a���Qn�k�2����,����n3(G'�#|���v*��Y˰��6.������i���b���
pȭ؅�k�:l����$�d��k�Lt�Y�4QOp0�������xH*���.��n�w��<�9�=���|�{�uZӦ*��-���<��S�I���cl8�Ͼ�)(�ܬʒ�[��������TVQEL��m'���I��������pouP�# �̈́5~��������L0�����*�%��sl�����0�dp���/{�)m���UXSs�)aA��y�ibA�v��J�^6���p�I���Y<�-
�K.�E�1�v� *o5a,�����)�ĵ�\*AلQ��ra�L������F�~N��� 3��R�DD]�6yPN~�6�0���G�����rJp��ꈁ]+����Fv��աd��I��_I&�i�У|
��%��֑��3J"�z�<�#?��/qs����_j
q�#V:"H忶�q��<Y��'qޱ6^-�r�6���R��;��DH֝�H��?����vYmm�r�_�w��>��|lc�;�ӋY Z{�̔�M�fV��?6�]�]����	�l.T�hُf�j��e��=P��O_o�W�`�i90V�s�	9d-�|5��,�	9W%=7�n{��M��)�˚&��y������[P���1v�B�1���PM��e� �X��z*��,�w]�U���3���0?���ft�x�����D��\#.L�r��i�U��(U�!��Z��ts��t�ٽ�4Dy�%���Y	 �TAy��K�v��B@IY,�zRY)�:�[_�q��N��m��垗��"Q�b��vY��?�,�^$e�JP��>| w���7��\Kz�9^ zE|2ه���c�SY��ђ-�����ZZ@8����^{��B(�,���"�~q[2 �@�R	#��}�u^ӏ�]�:��p��d���_+"7�<��1�,d]�O]<��IH�p"Ūa�j��d��a0�lFŊ��Ur�?4eY��?GX$%@hN�?��� ��'Sy�4��O��`/��%�_����?6_��4�K���e8nLVKE���