XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����u�����D�.2�0�\5����s�%��7�^�m�M�a2�C_W~,G�G/<�P��5.��(+S�*h������F�?-?S�ܱ�F�Q�q���<�,Y�I�����/�.�8F�KK8<�%
�&`�sNjА6�$��p�%�ioZȤ��|L��"�w�r��#�Ȃ��3��ްPW����A�����0Y���	_��X�h6�I2.��ܑV�u�8��<�z٧wE7�L?������,/J�����	���C:��#�?7ai-���t_��/�b[���Yj��?��˭W��cLj|X�`_���e�(�p���X`޶S������\�Kf*(GliJm��Z%��3}�3�A�Qwֻ�[��9r�\+1��/���e<�cEU�|:ui����m�+�U(�߃�ᚂ����l�����]v����Bn�Z"Ou��_�5�"��P=9-1?r����^]���sS�bY���G���r�
��T�N6!��Zz/f�˵0��G��*�660�0 ��u#�@���cr�W�I�gQ`+��.���n[{�~b b��ZIL�}�RF�t�a��W��礹��k9wYρ#���.���;Y�����V�8�+������Gvn��l7�o��Az����EJH��
H�$H_��ud� q��y�Z�f��c=ϰ$DnL��Z��^8W?��M��v�F4��@5m�A�=�Is��;�&��N���~�j�~���XlxVHYEB    a037    1fe0<�p���oX��d���C�cN�9��pR@���ۍ�w�f�w�qc���J�ª,��-�J���5ԅ�%�����I�	T|�� u҉�G-�����%���"��M��B����@Ԝ@G�E�X��EH%4)��}�����U�C���9�8eX��+@�0��	�u�VO�����1�aW�;��q����5׻{�����uUxxVkc�r�B؎�U�_4��'��J��m3\1?��7PAqL�*ڪ���ܩqo����^��>��^�Q�6-n"��E݅5�l�W��P^����9�p,���i�1�;i��Q�;~�GI@���_����n�۪� D�C� ���l��7�BD0gLZ��9*a1U����b�㷸��?p�SMs�d�>�fʷ��XD��s��w�8:�T��x�t�Z�Iv�hF��»��x#��J�z\��>�Y�a�S������<��'��� ��A rաؗ���d����O���q�V}��K��8_*t��Iқ�ָ���;�R���_�b,�v��v3�t|���g�|��%u���h��7ʞ�	A��pH��8z��H��*���6��F��*B�h�bD�<����7~@��6��\<�ʳ�k�>?��,T�s�i��:�W�]�>�� �u������'H�`��`�8�������ID�+qRy��|y���1Q��?�d�9J�d[Y������`9�be����s26_=L�;���t6�����٧�{t�X��v�Ե°��/1���)�rz6�}��m�ܘ���gdɬgq�86Kь����2���|��	��K��"J�K��o���H���
���%g���Cѹ�L���O�օ���U1ę	p�l%ry���NX�v�(��|�|�;[���  иDQ�p��g�ʯ����ӛ�h�I�(��k�I3�ƨ��r|���o�ׅ<'7�2�������fX�@d�g����q6na�b$5�FI��m#��MP|EBI������� �\{��Mʅ!�P�q\m�um�C�6�g���J�9��F�.�7{Iv�f���,]�i�-�!�v+G��ՌM�/�B�'-�:r����繮=^@tӥ<����Hio�_u�(�JT��< �h��� +������C�0L�
���aR߽Ľ�y~>d=AW�r�-+�ڰ�È{�L>����K5 ��O��W����"�@d�;��{Vp��ZX���*^Wֳ%�Yc,O���R)%��x��L� U��	r1)�
��`!�F�teY�c*D�~���'���PG�[)�Ջ�c�z�(U����rtB������`����\�Q������B�ʬY!v�U�l"(���e�~��n:�p��)��M��Gn,U�A�Rg���!�ZwL�h)��<�1��x�ȧ��Ct1�*2��ͺ��u鞏 ^'H�d�M��dN?�y&�b�B����ݪ��xY�,���n�5��#�-�ܕ�"����o#��P7إ>Gu��4���S ����r��`�a~X��AN�e[cS9�;p�J[�L5ә�?B>D�f����n��@4p>��x���i$���u�����F���������۰��:�h�ڀ�^x���JSOٔ!�#\{@����͝�Y����2�����}C䶌P��k�-�GZB�{3w̛�o♟����b)�cI"�ٷ��|�$������8W��*B�pU5Wi�Oi������-���qN[P �ps�XD����9�ݚ��m�b@2ި@	��L�X���������AS�(E+{��� �!�;Ol��4��\3��4�
a&���t�l���c;R��N���N]�k#�y)n�g��5���	b���1�c��;g�Ȱʝn8����d��i���A��Pd[ �m��K�@Ǫ�>�dt�E�m9�|������SD~%]��<܏pux�@� Û4�b���7J���,� N�$b�h���f�H>8 ��,��[f�h5P���M��4LZ����,?����#��x�j���[����0A���OS��U�|2ϫ���9��U��8��g������T�@ ���_�&�,�Gw٤�~��T�vf���S=,�)τ�3=���{�)ռ�ʓ}mCr���~�d � {]C��~�@�)4�+��/8��[zvn�c������9�,����T�Q`���&`9F�-�0K�o��|�+4�;G����iR�����3�o��ў^~E�%�l�q,��@���=�{
�g2���JcŐ�)q��l֣���r-�uټZ�:@��@�/y�O��-�vm/q|��QZC��~��@j?��6!��3�cy��!̐ �p���4n�@�;��jߵe=�^�ZT����I~��z��L�4��A{w��'��
9h	��3��F��NetI|~�[H$b��N��譫3z����������6��������w�K�
Ʌ�[r��q#�ӿ��M���{��1g���}��}��a�߇2��7w�=���nP\���r��L'W�)'������u���b�R�$�2m�(��4lC�| UF)~�{�<�cS�R�:�~�0$_H� ls˄��S?��$-�9��>��7��q}�Y�A��W�J��B�����0��?VAu7gLܣ"y*�m��F|7C�y���;��"�R�;q��2\����d�5�`��̧#�1��D�B3����-5k��o��֊��;R�S�;	\�MK�T���l�C�'-��^��p5�ދ�9����/1&��.��ֈ-_:l㢬��?�gX��>3O�R�U�&AS+��uG�*m����a����^���V&u�S���R��au�����O9(|d/fb�mg�5U�~�B��T�T�MM���f�9]���%X ���|�X���u�	��2
�?$B�����4Q*�鎭[��{����l9"C�J�# �;�s�a��}�;������$��'ѯ�;|&���MR+��������E�0��H09�) M0� 8	6V�!@+p{XS�@H��6�=�)rd<,���T�ݟK|�[�)��h�<��
�끃��kQ��*�9�z���ˤ* e؍��ł� ��UM�8���l��8w�'��Oc|�f���a�Y����6�c{FT���Z�q�W�u|��?�*83�~�[��M4�
MP}��p@iwL��}��r�d%��!
���M��\��ⴁ�i��Azg�2�f ���/��G02Tg����=dB\������}�q����(���4�CD.��r�L���I!-���OMׅ��eO�F4��:�Gj�$F@���p�<��s�KT��C���я)Ri/�ߕ�w�o����$��A� �Ih���rh�9�Þ|��Y�mDG���Ԭ���g~(�[���5(�KA�~�oD`s������䮐m0��d!B�ZkR�$U�|Jx����Ԅ��pX\[�]'U���v�k6*�D0��3�cWݦĈJ�����svH�Bۿ��^�m	�ʾ�45�V03��d_��:`m�`>�����4���eU��=�۲d� ��N�;����&<љ}�$�2K�-�81r��W�|O�-{,9������+��j��[�͛�X�#�CZ�Pi��Uo��|t�C�^3v�N��hQO�968�ԡ�K&a�����PST�w?п��z�,s�ь��(��J
�Я��iT����a��qwO��	k�K���_��w�ƕn�Σ8ĜU���bM��r�2��+V׷��T#U�M��Ky�ȣ8⶚�Ԏ��q�J�e�W�<��<�W�e�(1[�/C��o�$�(o�[�����-V}�@��VC+��X���=�A^�`QKE����q���§b� _t��+�޴�ԶV�s���v�m�-D+�x�C� �c6#�`�o�l��5��=�^A�^Ԣ2	v�}�'K���&#/9�|�ۅ>��0�7��Z6 _l��q��o���/]:CoYϪ�`��ָ������آ�AG�M�Ouu�J#Ƙ��2�����T���6�n��X���>�:�)+AHͮ
����e�VВ��)Ǔ8Cj)��~yU��4�#�C�{V��ͽ��S�<7=��ӫC�8�`��/��f���BY��<�-Ys�7��jp�O�$�\�PxZߩ�@�ED ��sk��P'r����?h�s�o�Nn�3^��D���w�R3Y��O���Y��y����@�m��(��щ��=6�J�! <�]%��*F6��#Q� Y� "jA���'v P��]}�o0���iE��5X͚K�7�чU�U�q	���=G0k�ч�}m�ߤh�H���(af[w�R8��^-�ӂ�r*�O�͍��H���y��h�G��m�����LCܙU���f��������ώ&�_l��rc}��0��>@ձEX&�`��nfb
����1X�N�x�5��!>J�h�����.ak�FɁ!�Kq�\16�� -��}��>x����-����2��>~���J��"G�{y��ӠT�μ�N!��D�V)���A�Ϭ��ɪ�g�2-��8�0�Q��Xne6Q�� ��J�.1D!_J�]e��A���)��Jj��g$����p�֮夬�u!�Ѣ�P�c�	:����7���}�V��w�G�K��^/8���5N�Cb����n� �����j����z+�h�/qTn�J~b@��-���~�Y�Ev�=��1�4m�^���������ġ~~�gK�"�:o"���]s�����+]��%�'��kʤS��,�1[��l}g����벵A�J�-vq����9�4�g�c�z v��H���\<�hd��w`ꌱ�:��!S3d8�%:!�S�6D
%��̀����z�.@�h�d�>�Ȧ�Í���VȾ�n�f�|q�X��e��IemfJ��!gg?�~�]�'9�'j�����SW�/3{�yl��0��}����U*o}G^"N�2ցޑw7���m�n�p*��6M8�+�Ì����2�����g����V+9��Ɵd�7��߅;KC�ۋ��Hb�	Q��2�����Bznќ�����N������]�S�KbmʰӋ���Bi ��J��>� �����B�6�PY����N�b�/^ًWR
H2�]�
�Q�VyH�e��:�DdkgO-|��]��l�)b����z��!��
���y�y@���Z�l�v�;�w��bt{�>b�V���(����4����-�Z��2{�"=*x���4�r�q�tm�H�1F��~��͜�0d��~,�r��庖G��u�U�?�bp��`wt�Y��Z]m�+_ۃ� _!�������_YeK���--T�����\� 2�ɧĕ-'��L�d5���YE��Knm���Һ�|��_#%�p�8˸�Ku��ݓ����,�#��]�$�L/�Ok��w1p

�V��$���N*D���w�����A�V���P��QF��?:�(�n��Xן���Ʈ[��p�~��G��#=-�ƪ��xg�#��+Ʒ�rX���`�2�ɾ�+��Ė)pɪW�%�!s\�ݣOΩ�}��W1r���s���j�������G,Ս��sx(���:d�L��vG�F3�.��w�0����W(eS���O%[��&��E�<Ƚ^�m��R�k$'�?#�O�ޜ�W�.v�Q���WI@WB�},��,�y0�ˬk��vA0�����7�-y�� t?�� o���ߨwchz@���u⪿�"3�J�Z?��'g3?�����L�f�ɳ{J
ᥩqkX����@��kM���ǐ��ྑ��6�dA6���I���-�LzZ�]T�[�r�Z��a�u(�A�2����=� ��> ){���ÊSi�{|N�o��SÇ�l[G�V�J}=:Ƕ	��4���w���e)"1���0����e:���B9��q[�k~c�0&���o���R7��U�f)�e �#ܿ�ŷ���O$�l7c�<�����#�/��7._\Ј@p
������j4b���t˕h�I8����T3�(�]�N�.�rJ1��%&�������%��9��.������d�XS.�^~��KϐP��t��v+��yBNlq�Co��?Q���)�H2n6v�+�@��A3v]~P5Y��t�tB�-|�A����5_��J>�fTw�����;�6����beS�P�DΒF�
��Ş�1�NAf�+�8�K�̸l����}n�C,wn~g��Bf؂���'h���z�	�o�)�`Z�/!�-��?�V�]$��Y��~�G���i�3�ܲ�}� ���)#T��צL���#*�lO|U��X��g����c.�К�4��2�9Y._��6����5|+K����09|V�PóP��r�o�;�`t?T�� �ea����1:�me�"���k��X�Q�3���h}e�$%�^�e��faY�	gH�%JvE�F%>TO0V�d�Bf�D�Ť];�frۺ�J�uZ�i��U�K�ԕu�2�"��>Q�� Q��e�R���I�~���i6X��]����4�su��	���N�j>U��������({���	%�+�_j�u�w�粛�{�U�䳘�}���`�Ъ�j�.�?��1W�Cg�fn�
�.P���X\��8�%`dh�k��G�{a:�e���߸���^�L��0<�� ~S��JC�&�����8���A��9�2��ʥ�#�O�#�y
4�m��PtC>r�[����/+H�Y-���$x��oD�㴺��`������(͜k>����M���q��f����U����4�wZr�f��i��`���Yk�ae���~��<R�����+K@���w4�Vf)"D�Oa����6��உ\'��`��>)G�K��i��osԚ�bE��sz[�q��6FG��{�������v���ʂ��3��u��v{��j4Pa�*���;=��he\��u�hܝM��<ie}6z�����$��FB��
�	T�$�F�_�-3�������I;�n�/'����%�F��(|L3�U��,^q]��C�m&������# |R�$� xw�E����=m�	���.wZb���u�w����hj4G��W�D��UOz�K�@�:G�R��YyV�;|�?�6ۮ�Kj����I1�NQ-��h���[�1����8fG��&�_c��v��&= ��P1���`U��Nz'��[�@[�'l�����R͓\� 8�Wj�{�\���-އ�c����8^��+6[��I��_!�EG���Þu���c�������CVpz��ouXE|l�)/��O �Z<rz~��3y븷�4,��u��q�9v�뚯I��U�95BO��2�p"��_v%4Z�u�v����آd�z���G���^׉*tk�"�A �v�6���.N#�g���X��|c�Q�K fW!�n�a�v0,ZjTL��p��J4p�+�Z��Oo��������C̊%�&4��u\	 5s���r�ٱear�v/m���.d��� ک}.�Y��[��y�����j��)���z�`xȥ�T�ɶe���=2V���O�Qy�*�<���c��rH7/;BC(��Q�DQ2�_[��������Lh�H���h�r�*l�W@\���Yr\��GZ4�)�K�(wf�?���;K���GĲ�里�A�G�$'2�kl����`�e`͗Z,������x-G��L�	3E���
�@򊘴�Ug�B��N���������#���Z#Z#��^�7�p�2}pd�5ɀ^�X�O!�w_�rd! �S?�I��`��땨�@ŭ8p��G�5K}�ŗY3fh�gvHA�M���u\�+�M��O%n��� �@ӯ�GL�I�r2��We�_f�L�U�����ڿ�	��M�