XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��H�b�͆��آD"��^��yJ��q�� �id���D;�+�C��\j����`�@�3+��<�������Dn�I�~�msU��$b"��E#�n�l<5���V��_�8a���B~l�r��R�l}bQLI@���Y~2��.$�
o��n��&�$����\����y������z���u�A+cfLH�t��vR�L�W�:~!� ��/��39�_�S7zb)��Q�x7�r\��3/�8(8c�"�I̊����L�+]�J�u������6���zs[����#xb0̄~H6=c0�G,l&�$�<q�Cy�W����D��M�6[Z4�f�c���R��>z��1qN.I���Kw�{)T���_K;�b~l��ә1���=
0�g�2
*+x�lx��%�M�Ta� �/Z��4�]RB߬q���������J�g�����)eLJDK��ʂ2�pj�,���A���r�(-��9�m����I��2����m��Ck��꯹�p�b۱R���ue��Q9�Yٻ��u��j��^ʢ�L�q�8�f��\a��_n���/�cQ�f�zh�9�[�6;N%ir���⩎@���`���'5�'�yĶQ/��ͱ�z>qΌ�德�#��If�҄2w;�2 �m�)�z*�g,�Uܐ��dlV�$PԚ�|�Y��+�׺�2!ͪ�<P�Xq`#f�A�yQ� �l*��:�o�9Ϸ��Hh5�t����Y��-�o'( ���-�l�V�fXlxVHYEB    95d3    18d0��=���;o�i���	���?�'�����4g�I�XXH"�t���bg���1hQq#�v���q u�(P��Ō�@��2ff�Z���4�(��%����	�V8�f��ˍ�\�A��	�p���Z6�ԩi�Q~w״���&l:&���6)�J�'��j���~|S_�gN��73�*��cT:������x�7�0Ƥ�,J�a~[�RB�����[, �x/N:��v�T*�.�@Ԧ��g�E��rZ�<o���8�Q�w�} [�T��;���9��a�U��l�������Sc!��$S�Sd�K�IM<C��2�,
���-���;�ho���Θ>n�x�?��,�>>+�Մ�S��}Xt�y�l`��&��prm����1?J��<x>�%�� *��"2��K��:���:�%���� *Q��zH�?�F���u�n�1G�4QY�'w�{��kp
PaYk0ғ�[0���S6�9r�4qy:�c�F`��P��"z��l�M�T,��������B���]�z�:��+�p��7�P��	,ǜ��>n�h����<�A��}��Ȩ	�5�x���0a��`V��5�Δn�C&��^�ev^
��순�w`���Ƥ)��%Pi&�q|>�U�u��3$)ۀ`I( n�R���>+.��~XY�;|d��@�����	� |2�k��b��!��ڮ���κRd"��ڂ6���N�
s���Jy6~���lZ#�s�ަ)i��)�0o+E���e�-������ �;8xz��o`*2�F�-�F�6��Q�4/*ȇ#x�����h�o�-�������^Q�7�����=�Qݪ%j�"�$����sX�T�G�
k�YA�U�Pҡ��_�dAQ�5��ϰV-����&�{��!�d��Y�u��E�뫺���z��߲ARh��^?*h�eC�)�FG�d��Oquy�_;�c?x�r��_ ���8���d֐Ħ�A�WQ6�/u��c����\����0�'�[O�B�4%`q�����:�L~GVm���3�p�%�%��\%U�9�=��[�J�f4`u��h�+�/�7f
�-}Jc:�,�0�mԃ�J����5) ��3MH�����tɒN�26V��Θ#hlT �S�v�=��nǜ�K\��cH̷��'��SBh��'�غu����5�a#�����R���%^��dگ���8�.�U�6l��i$D�70���`B�i�Bq=f�P�ό��6�_s��-�gR�Ec�d��؇8釃My��:sN��='��~M")C��&Ls�O	�%��N�Ycs��FZ��|�XH �Q�x�)'�e���g�Q�� �i�7�~���~)ښ@9]�<�e-r~�m���8��IsM&mr�'S���l�وr�l\fA�(-��hh'C��f�����`RPΤjP���&6 ���I����(�*f'��Y��n������lm���؊�qv%?�	�<*X�$�v!J5Nh��%/����m <x�փ(�󿽩 ���j(��i�"���� e�"O���C�b[�	i�\
�A動>�R~��_�i��`g��\�>"���!�VB]?/=JW�������_�1U/���*�CН������Z��[Ԕ��F�+��2s�<�mʁbNܨ��,��Ś�$l����Ls�G��.��5O�:�%���P�F�]X��f��1����B�~���S
�X<��$����]4! ogQ�I��k�/��	�Б����-r)?�}�}H(�H��j[!ќJ�G=p�e��8�G��9&�K�n��r�y�x(�x�gS�J�T]@܆��R�m��f^@����B��}9�Mg:����L4Ŝ<F�{~�tE�
��3:|ǺN��g�����[�����v���:5�R�Z�^�®S���=����d4�=Ux;5���˼{��jF\�:�	�J<j��w�C���Hd{�k��Im�۩|T���yr���d�xu�2v�z�co&�-	J��i6��fQ�>R�X�"`�	�/��7��|/�U����ܨ
e敓��'k��P��&�c��H�MV���+u��ja0f��
��J\]�}^����%�vR�O)�
gC`��Ü��;���k�J'x�b���^~���"�]�U:�f�ޭ�p.mC������֋J'��N��vt���e~BQ�V�M����_:w�3_95,'O�vO3-*�]J�����[���i\�SS<���bØ=���fKpdgy�%�hz�g������W�ⶾ	�P�79��I^�>��8���x��/�OA�=v��W4�0�P�<��t,�ӭ�i�@�dv��c&�*J_9N.>��ӥ7�@E��Zv����
���VAO�\+zK���:¶+g����cHY���!��a$Yil]�m�'�?�B��N�����0�A:9mK�O��ȷ2��+�6��R�[N)�X2h�����AĤyں�*>�Wn��_쌗�}ƶ^�Cm����~��ʹ0]}��U^#�:��KEB����2�[<-�Ů�\X7�w_F��"ԛ�Q�*zI:iT�40�Ҿ'�ꎺ[y��-ԋShg��l:���r�"��+�QZGR�ŭ��]݇�=E�B8��6S�])�d�w�"z�� ޲tP�լ��j繟�_b�`��ld�1j�o�0�C�2�+�E���*�]��~�]A���]@��gƃt#��0!w�&N�e��BU���樓T3��n>�E8���>6^ �v�4àՔ����Z@���7�+�=U��P�Kao:��[�-��L�a��j|'�8#�	x��Ĉg�%I�Y�k�9K9>�5��!W����֋�c��dg��R��.��X��@E�4�~�$א2T%�Cb�p��.A4V�ê�́��@��_"0yN��<���C�$��a=zQzg��q#�& �Z���A3rs�I/ڦS	zMlN�V:�Hu09���L f7Z�͵#Ȯ��Ѣ�8td�W�QJ�l,5n2��U��8�\s�I�my�(�"���zӖ�'��F�
.�<��L��7�v�ݞ=�V�FW�0ʧ�{���hM ��J��
<�4��\,���&7ŧ��x�؏���߆��6���U�J���x�������'�#%���4�rl�8���$#l��b􎄐�3M� _~�^�3*�|o�Վ��X)�p�8'3����k��LbfS[�_x�a�M�c߉H���P�'5ѧ��7u���d�6Ee��{�&z���
��4�	r�Y/IH�v���0�ͬ�^m�5}�_M.fe��Iks��� �-1��v
Op�)��z���w��-K�d�ދ}0�I��{G��~4*��G#.8�4��2=��ԫbd�u3��3�\��x�����h�K�I:�(A��q�=39��k3
��p�1�\xs
ϋ|��h���%̙�`$�c�)��|�f�,�&���-$R����Q����&�:��﫴�3�䲍�����)7~��x�vt�!cs�L'�_6��������� �'���0�F¶Mfw�}���a bq�,:n6��.>Rv�n><�n�g4���OF���� ,�2���%��jv���ײ�>���t�i�0>tڔ?�,l��cZ׵.�ˎ���O��2mԏ���:�,��Vӣb�n(���A���)�;&ݽ��=�>�ZaE�71�Sh��<Bm�Q>/�_u�x��D2_��40�:������ߥ��f������	�L�GrM�r�a�6*
�\�a��x�ֵ~��۶*(��H?�x�r�Zg� 1g�/�S��`��;��l��/`�t�io��B26|��.���q�ِ���L�(�m��F�����M>�/�jf�Pꈀ9����WW�`�|@�R9s��F�0,Y�Wo�k�Nw �=i��~�`zI\2�>�/�3.w-U����Z?��ޖ>�}�h��/I�K��RoE����L�+��yؿ���
m��=���&�o��j��G�5"�?W���2aW0�)"����~���y:�
K�6}"�s� xn�]�{&6����Nx�O��2��H�lG� @.G���V)��6�yb�zy)q�UP��h=\���k&H���j��İoD��t��=�#!�!�1�����Gǿ�p7#2�%����7g�O��t���ұ��.̓��q�~�}�^U�6bE�x�A���D��)�J:	<Y�\u(�?+ȁ�J��d�����k�A2KZ��>*JXZ�X��F�6�h�$"i�>=�n-K��� �="B;Wq���G���Ǣ�t�������_��k�{!Y���t��P��G���R��P��&D[�*���~�����N���U&��z�-N�e�/�aQę��jΌ"}���>G=r%�9�l2QÕ��9��2aŁ���%q~��i�~6���z��`f�*�횷4�oV\˯'�G��R�G����7n��Q%b]:���t���x�fri��ZP���Hf�nُ�d.��L� �����Y�<|��D7��4֞K��r����ކ� �z`�iH��%�w5�ԬwH�~���7��r丙Z����ܡLY�n%[�����>����q���E�i���z��ύ�=��83�.)�]gSP�mθH"*ЮvG�=�*ȏ�BN��%�Ε�tI<b+�1�����xtW�ˍ�6�x��ۋZGN`�����B�a�N*�ґ�佾A�o/�g�o����g�k|�_���%p�R{1r[��z�}����Ⱦo�2�W*��_�LNV~��3��)l���uFT�a98�C�B۶l�����53�V�Άo`|{L�k���Xu�� E(�.a�/��P�����
[�qc���:�$�5[�i�J�OقS����@s�������aT�V`��I�4��o�ͥC�B����9���1��i��/T3!j�SҚ3�Юal�!B�?��_�x�V��'�+�(��V�vot�~�[�1�r"��c븻+��>��86�����z"$b?�j�#�h�қp���
�I�!P��$�o�[�k���(ێ���e�]X���z�9��U�Bos�����������c蔴�w���f�$]_�[�~��Wiа�d�s	g\�õ:;�����CL�L�o� �2�Ւ�_��6�J�!��n*�"f��W����S�\�cQ>�}����׮�Ҳ�1��*�܋�/��/|�?`~JI�;+.�Wt�@9��cS"mcb�G�ht�%k���ꔇߚǢ�HV{�!	�ѐ��#6�[��罤c��΀$��ˮ�0�s��V�,�}2{{E�x��E�=���i��'ԧm^we%�;�� ]N�����+�m����ͫ���w��4�l�z`�V�O��Cf�S�	�.�#�?~�����N�
�?��qĥO!��{,D�U�55
��~S��1n�Jݬ4�^ª�C}�T�<PJ�䛱2�Ӭu4�<2��N�%d�0}��S"be��n]�j=��Z�b�=�����^A�@&R���0���[8�<�d��l�h�D������b����2ǲK�e���v屍E�؛@����ȶY��\����j��F.Y�r�h��p� ��\�4G4)�LD�%4�h���_�p�̹���GE����gx��A��s�G���H��}��NӋ��Mի�C1%<H#u��ySlF�����s�[�A�"�-��TŚ9%�}��׉��;ұ�W�K@9��yo�B�&�IW�6�{�D4���NM�#�J�S�|'�' ��������S���؎��#A��%�E�7L!���,'v;��]xg:7`�?�,���w����^�b�;J7X'�𥘽.
��3H2&q(�t[�e�E
��R�i�4bn�0#���7ޟ������Ѡ_�&_������=����G�q�NI����&��}���\b����-�kqA�����6*M4���s_"a()ˢ6��i�����f�7���� +�w���TK�SU�]j�
\�K*%r&�~I�E	F�ٹj+8�s���8�\=h�Q��~�������#J�n��0uT��px��>�޿#��?J��h��}��ڂs]�6灩����E�mow$v"J��>�S�&��'e]}o�h� &���7�Nj�	���`���F͠����ճRƷ�2���2�S��0���NT �f�T�%�߷�	y�|�w0����Dv_S��,��e�iV�c�SYv����
j)c"�f��