XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v�\T�A]�-߈�|��r��$��%ܳ����O�˶?�m��)�k��Ae,���8w��e_��]�煠�����B[�����j8��e��D�<�W���uر@�_S���A�x_�[�]X�ōm�w��wB��LD:Lבy����Ȫ�y'z [�B�xƏR�|�������B�?�41f���u��zi�{�{�x��لp�d%��[>��b"�<_ّcN>���%L8�6�5�0�d!	��?/zD���@��=�M�BX5�Y�@��+�-���_dSl���-���Z|�⻤/��^CMS��g ��Ќ��*oGQ��R�-���5X"��}� �Q��jX�n��
˅TYd��I�F���B)�̙7�����mN\$60���DF�MW�.|�.��
L>Yg�:��Ja�/�	4�N
[��S�������K4���?ĩ�v��9��v����s�0������Z���.;4�G)M��UW@����z&Ԙ\7|�
n���i�����L=�zE�t�P"��N�ݘ�׭4w%
Bᤸ�/	��gZ��d�y��)5�quU�Ŧ:v��e)To��,�!�A��m�+T\��v��R�Iԅr�1�/�6��RV�Cb�Y`�m)�����G �E��mE�U��E4����:��2���[�ϩ�����ܽU N/S����h���8Y�k6EI!Wz�"��C�f�R)�����'E��"����L-�W�Q��� �a�=vKx�A�ڥ+%�XlxVHYEB    fa00    2040n�\C�Q<��%��|�NO8n�z*�X+з��W�7E谥��sδ4�\���C������+	����wM�!��SƊ��LHv^���r^�����)�Y��;��q�T����R�v�|ǒ��Z�ϰ�[Prl�0�ɜ1V����ֲ�c�?;6��)!�N���xG�zU�֛����.�c1+]�h���Ѽ�J�s��_�2�k���O�al&�s��*67�vT��l'�Ȃb���
QѼo��a#�tyr��]X 7l����E͆
E�
�� ���^s£��J��ĊKJ��9t@҄sn�u����o����$/�Z�km���%¼��D/6 s�p��]Q�n��D� x��QcEGߝ�I�� X��UA[_��q������4����UjU�?��PB��/y�!{A�3��Z�~�|��s(��:���Q�-V�Z���ñ�3B7A���������EV��¡�J��B�KH�}#�!���\3�Kp�a�����I��6H�s���Gt�k~O�.�V���ʺ&�? =.I��D� �Ƽ
�!j��I�Ry�C[]���b�9�	4��W�3U�[�@ڔ���3��g㲲��$s�U�0ގ	@�G��h�vD�fr�/�1��xg�F<���iݹ��i���V��Z���%E��^�I�Ñʐ,��_<�T�U�?�du6u���]�����o6ã����*�=NSC����.t�9ӧ�Ki�EX�$E�}!�LӪaG���p����x���@gD�׉L�NM�CoX}���/{��	������`�͌�����w����W�V�D���)��R�`�'��(�>����3i܎؅�z��Т�:Ҟ�e_{V�9+��f�'�ZB`Ɣ�y��fPbQJ���.2��w�0�T����y��Eݤ3:��=F�s�j����D{%�׃>h��|ЦТc�Z�d��7b]�3ʚ��I�:֞A���}�F��DwL�
���5���:[g��ӓ�����q��5�C�8L�b6���L�Ѧ�%�SHD�J��MY,&��9��:�
LM�
�/:�v��yt�ʓ쟟WXu!��)v#���>`���GUl���2��΄�W0��(����j��ʈ$I���ͮ�[�$�v�px`(�Uu+*��j�/�9�S�^4�Z��� �훸�mH�OE����l�8����%n�<������aFhf�ki�\��_����� �o�(6�Ř�i)q���_�GT,Ҧ�x��cT,�{���Dشg�}�	u�C���l����Q
X0X�ܦ���	�HX�1k��5G�j����9O2���b�ꇶ��ْ� z�K��0��(%���‧���:M�E+�r[�X��C�'CA-��\:&��w��n�0!�YC;2����<��[�otb{q��ݞ#�#�NnCe_��i�;aR���-���*�@���켼v۠��D�	{��|��ݝQz��i�4���˃��e�A���}K��=m"�&
	O Q/$߲Z+Ñ�>YB5���E��,�|���X߃�+���df���Rl-�_�)����|zn�v�5\�up�{����ٖ�$�1,���Z�-+��Z�!9͆���Ed�i��/>�Zv6�.�x���m�\�^u����|�����|=�ajU0d���
�$�*�x<���0����h�R��2,l�P�!�̱352����G{5 
وv��� �ёv����#(���_�:``8������-G7z�2�z-J�O�f|w�QC@�cG�q�4��ԥ-L���N�W�����hF��x�Y��4
~��y8��91��/�8+i����fĎ�L�7*�X�`��"���q��	^���K
�L ��xNSd�?�ٱH��#�Y�p��H�Y��Ù;��I���;�_�v3w�����Y6L����]�]�?�Q\C/����,�rKP��ӌ�  ���|�PT��^�m�i>��[�����h����cF?�O����7�YNn��������f�t��s3�&�����L^�_���j�'tg+}O4O>H1F���?R���붷�[�V(w�n�|���Ч�U���>��L�;�O���	�x��v�M;�6>�D��T��l1bI	��/W����;�~��'?5��H�x��>�L���"�����,ı�6=�� (P���T�B5�!b×w�y6#�s�>wHW�#�D9�%�@��Z\/e���Z�=��	u{+����o
����eɣ�s8������	d��K��+"�L���un���bG�*���'j�)X;!	�n,��'7����쾙�|�+'���b8�� �1��y�`4!%	7nVܹ��y(��P����)ћ��s�t�x�5��G;/���wՆ���L7���sh���#>��qBd`�1�b3VoM�aV��v�`vp���W9��x��v؜p�j ��G��' ��ۅ��D*�K��j�&�z]�jn�@���ʝU�	,��"�Π"7�Kj�g�Lв��Ӈ}�\�G�ɫ؛��ɞ,+Lx���at���ɯ����1#���Oaq9�q�\>y�D�9�\�tZ��Hp�G'�_W�n�ei��T
_?SS±����>�i���el%X K37��?�dU>My��f<��Ոb\IV�1�P�s�ă.B��_{q�/m0!,D՝/��K��Mөe��u�i���;u�P�8�2��xi���I�6�w9��e���Ye�4�S�h�`R	�g*���4�<�E����Wc�(��4$:�݂����];o:�W�07�w��u�^�&ǹP��Ŏ+h���-9T + ��8�*�O�	fQ�MM�w�s��W�������>�F�|�#��۶���	�B#��9�D�SN�����&y�cw?1t�a18@
Ĉ6;�ޠd[Ӫ4����*ח��8�]�*5�攢M��k�1���j�6	s�7"�w�L����/a�[��U��i�H9�n>��孛&T<�7�.���t�꺴К&:��gd�P��K���W����.4!��1�6+&2"�%k�F]�/��s���	~�����c�Dr���o�k�hP���+��	����͈7q*벣�$�L���F�E�SJ4�\��lF[�4��Zo���]�c"ށ��,��l���C����-��t�Ȟ�LE�������������"�$�xr��ґ�P:����#,�్ً�շ�Ys�|�Mq���s�<�-m��J��2g���E�L�H��:��09�:���U�ҝ+ϰ6
�~.�Mb1��ok��?
�'�f��}ص����X�{L��%�q��I�y�Ic-B��v�ܚR8�ʖ�!��:��Ss��
���w�����FYف���k�M�:��L��BFY�L4�J��=�[^�Sz�AEyKoWܦ7���*��t�H�D@�%���}�/�"���l�8�BQ�|���b��},sf�媯����3�KԢ	N��R�O�\�-�&':�V�QۉU�缱E0���+�|0��X�&����"Z /䨅�u�Sz%L�F��0��
e�:��š�p)���C��c�Q9;Ż[`)'A/T�+�JhzA+J�`Raw�[:���P��ߢ��y�����@\A�z�&�ʟ�o��e�q*E^_Ci�8��zF�������j48t��7mIx��V���� !\����o����Y��D׺~�ew����'Hz�"��������)��!�WR\�֢�;Xw���Y�+H�]�	�D�	U������7�t9�я�zH&�^دX��e�hx��C)06b3��^��-6�O7s/��B5G���˫+k';��bP��~2GI[铅�����E0��נCF���53��v fГ^0^�D3?��.�@Ʒ��C�w;�����M�w�|�-ɢ��s<���=�%QŲ�\��G��ahu`�����UF������N@ت��al�{c�4��g��{'�Z�.v����h�����A�����Д�(4����oj�~rJ��Ew[��)�$�����O�.I����`[��K��qMV�wVI�e"(A(tHyT�7K5\M�L'�ü��%^�ɛ��o���?LzZ���E{�7���0,�m�;�B��3�h;�����vW����\�;��N�U�T��0Ĉ�:���N�ͭ ��c�tޏ����O�6j�jF�c���@�z��y�	�Z�&
����8�]���W���&�݀�ʿ{j�-8����TF��7���4y�+ 	��,G�+�S�[����-�j�����5�rY$���+7��ϐ���R�H) >��?�� ���X�9ni��$(j�:�*��`��A���_���nקd�&e��[�2��+.���H�(�5�Y��h +���:n� �i��c�A�@Ȑu����\��I]���3a�AV�r�,`]QZ�m�A��t:��UX��R޹c���.I Yζl12�n$��˽x���`͉�����сf�݋)/���?�0w>�&[N�KΓk��^M���Z�E,����M���h�]Z��P� ������Zd)���&�ZP)X�kQ/���=3�>O2p����f��t�����H��<R@�f5>�u]5���f��> s�ʰ5��A�8�~���� ���.�^��EM:�&j8�T�����0����س<�_60I�Ph�!B�(̉�09ʿW%�SD�[��B���07�h��Ro���^���e8��s�����+���H��N3?ۀh�\BOuf^�9�A�}�+�~¥#��g���FÂ?8ur!xhb��}mffL]�Zє�z�e��D�\B����Ñ��cx����)WJ��ŀtOZ�n��`C\��"����iE����F1@W���Y~7��Z�4ِ������!{��H@R�3�)��n4�x�j�b��Zri ���G�F�m��� ��T������z�\Mvs�xK��uA+���	���z(�T�*�IU���T���sn�+ji{9[F�l4��#h�Ŧ��n'�o���<��P �<�M�0��i,��DI%�]q!*�"�9���O�"Tc5�d%�Aƒ��hd]a"e��.��*�q�ih�Q�bh�!z�B�ĭ�FhԻ+8$Q�����5н�1�ÿifq�qTy30�\��5=�\��ʱ<S�L8�%�K�"��(�_�	����l,?^�Q�+ٸތH�s���׊�b��)����vF96唝WgV:m\�]=Swv�=��!^�g38_{g�h�d��m��\T�Ne��)sɉ���B�.R$?���0o���Ŋ�;ZW��Ė�d�z�L���<ߺ@�����9�d�D�,�b�\��,��Rm`�;�I�����=�
�'�,�L��U���I1r1q���������F%��,4�NR|��S,�?�tA�cp�b�����I���!���-�
�~۴(����N�܊�pn�3�3\u��>s{�N��On�jp�/f���<}�����)����\@�� %�s�{e�F�0i�%=�)������=;�'�������Q����(�P�נױH�L&�j��������T�IL��c{�ّT˽3�J�Y��iq	f��Grvk�#�NU�tC��`1}�/�r�|:�e�<(�n !�x�8�F���ө�Rf��L���+0�k�o&+�h�	��f`r�s�!���+ϴ�+�� �yЋ��K�Z�% |wh���WbҒ��I�a/A�����/��A�yh��v�=��DF����!;�Ѵy7_�L��<M�1��ګ9@�����R�=��Y��U�HT��D����p
�������N��c�L��0�%��N�k�C�=Ozh3�A�c�
A�ϟ*���K�a<�ǉ��!�w��0<�G4�"Wa� �\�5��ci��n�PO0 ڴ6�z��]��nE�W7��Uv4Ge"�AR��׾>/�ߨ�/ Ba��Q�Jǒ�+�v�Z&)�d����!��#�&�#@M&� �[�)�]ʻO��!�����o�$Gd=F�e�%���ګd�C:ֺ��Ro��$�!g ���{Oo@q���9��զ\�X\5d�dڙpE�w_~�8/�3���T�,�]4�`d�$�!��rUU)�#�Z��a�m�
������x\C"�ᵨp��)��>L���*�k�SEM`��C�"L/�$�`��Z���r��(%6/�}_H�_=֡zr��z���W��]�O�8�ki�=�!p��R5j8B1�m;+SX�6b3�i��c�6��/���~��^g�"��L����H�H�{hףc�㥛PH������e<���i��:�i��K}'�*H�S�ґ=�#�� ��������s��E�����_.{����n���h8�4��E����=�Nڥ���2�
��<�m���39�[Q�ƛ}@P<7gO5p;	^j")��XC�?�x~TkS��l	[j�\]u؋bPLA�)Y��]!t��ʏv��W3�`cݴKG���Z��`Cd̡���*&���B�awV��/�AC̍�B���!B]����t��q�.v�E�L�`����jо��`�vť6�{�v�K�9��c��đ
�,�#.D7#`2�JWE�Dt�Pn��l�a�ٶv��?��8~@�Y�F쭕�B��î��q�8���`i�"^2��Ɲ4u萢�l�	�l>wn��k�˝�tnK��P�e�9i��/��Rf ��*q�7GԽr6��.ɧp���oGx�<]�E����?v9���Yk.�����?����rl
��̸"{�<W�q �`��#
�)�r�6��㻕u�%�]Xv�ܚ���(~��c���z9�@��w����=k����3r�rt+�_%��_P�ԟ��qAvJ���p����Z	~s�D�ȉ������.�Ǡ���l���F〿L�aB��jm\�]��ޠ'�Ycx3������/�j��I�S�N���P��1��9W�H:(�4x	������{{�XXl�� �0	�8<ۋ����v��"(kq$h���e|�'I�VìKx���<��a�f��Wy���=W2{�����G��
=�B;�O�D���������)���N���k�S�?F�S�(v��;PiE����ON2�?�$���M�{�{��X��l�
���v�r>�	�*���+@�$��QR2��
PAs��]�^� �;�������mʯ�(l��,(��Ul�>C"Ǌ*�С�X�k8�P������%� �A{l���%��Sg������N�61NyKbT�$P�r.j��6Hi�[����<c!�Cs7>� �fI���`��!%,�uL���433����!�	��
�*�HOM�պ��u���>u�X�|���RH/��	Ӷs{� �W�N�����㜯�>�7�;4�u��{�o��`i[��x��O��*�3'�A*aŐ��������t��z����Iz�Yf4�2�Giw�\����㍜4;��ほZ�4�81����Hj �¶��kQW cĹ��#-A��� ��{�ij�Ӹ��|��^У+W�C��b~K|���o�f�ɫ�ࡖ���eY �}���fk��e��ё'XM/.GG� 
Cb��<uG��ċ�iYi��e�"l����{PT����,"�A�A|�o��C����
����z��7p���4j@�!�����=L�zm6PNl��k�*7�	Vi�UsX�?T[gP!���&��ҞǴQO��VLUU»�����a�Z���%ēr� 4���ga��H�^��[L�B����#�ic*x͑mB�_n�_�z��B�TS�\u��Iw/������b�ָZ�>��ژ��c�>X�F�tvp��?Rɺ��ZJ���p�Ih��<���\��m����%.[]�]�iR��Bt��|���1�ܗpD�ż��vE@&It��TW#:
��Ս�f�<b�(�i��Z��6#�ѷ�/,r&�f
��}��Fx�[1���y ,�״�[KA���&d¶X*E��̿��/��ԮiO[�"φY~ K͇� �R�XlxVHYEB    4f62     b50��uY�����?��0�Hh܂�=qyZ�IAF{����c֏�~|��7���O獓L1B[��-�\��#U�1W�2XU�u�j&^ �cmL��UGs�~/9/�w=|�Tc˻���PMjhôbRH����T(�Z�k�:�\+�M6z,NBZ�������/���%w 	���*��;٢���e��\R�������&RTXN�ԇJ�q�N���釘x��V��\�L�
����Ֆ��A�2��=����I,�u}�"�H����%]�P�~�iGQN6zJ:p�3s�O��0c�7ᆔ/*�@ݰ���yMf����;���л�l��K�	ID�%?�:�����k�ޜ!>2W{��t��!�8ߜ��c�����a���#��~���z��,��ҭ��?c��)2���I�H�|���!��?
�%'�B�=�BVKͳ�+ՁwF�r�LV"�U�u6�2Eu���]�~1A�wZ-E�@�f��q�ʣo�^nة��`+���{(_b���.�\nO�2�ל\#�AzC��H��;�]Zd�M���`YhOg��Ϯ���W�:R�K��5jм����c��;��mI�e�=~IA�N1��������iT�T�.���k��-���/��XjzYD��G��S	0.��+���@2uͫɀ�#�uv�~��`���3wد��Y=����1d@
<�ҶXs�du�S&��I�VPMZh`[d4[4�I!��#������Fh��V`�_��hLh��˷:� ��x���Ee�P�⥥F�s�«5�����U"��s-+C9񌦻�\)x�o��&�x�K"*��CE8A1Ƙ��T�rڶ��W���A�;�^� 	���1SWMW�4"
��V�&ڸ�ӎ�9F�D���FAv=HG� L�o�=Z����R^7y�/�p�SQE�Eڔ�LI�ka��
Ȅ50�k�B�dƴU W�>t7�_���E�#�2��q"����pZ�\L<�6�����@��=w����Os(����q��3��v���k0Ç eD��&T7z�C�P�S{ɇ.	޸�V���w lP��o&@UZ2�_J^��)����ehx�lM�ql�ӫʑ�^x2�p�8��y�g�W 
�r�<�Q*.�5M2��-Ε�!�t��g<MQF�s[��Ć�2qO�q*�v��}��f+�Ax�Xc~�>+�19�O���)s�/�9��~5h��2r�pl8��B��j#����B�fY�H���/��F%������"�{>���a��1Q�����~X��X�ŵVW�����Q�!^2|Չ���^W꿗F�2�wċrl��.��sU����lqC3T}[x����L���`��"g�A�ub���=�����N�����R`ι9y��s� �@�2翓�M�/������3����̧����t	ڵ*;����U������wdN���˄#�o��˭N�Vȹz{������^�w�i��DR�y2�M��}�]&��PH�x��
R�Y���u0��i�`6�2קÊ"�c�Y��w�ؗQ����\���� ˲��>�nɡ�j�Z����C��C.��*#�PJ�d�8�MO
�����K�V)/�T�����kg�GD	t7�Y W-��'ڌ�ďԺY�ǵ��ߔ��9Dh�,}��XR�nӅ�+Ƞ)4�`��'g���)��rr� az�r�ǒY)����;��@4Վ�t������� �v���]��s@��U<�Z'��)�8����`�c�TD%Řç���Uzw��7�o�B�>����Kx���U6����˗�>���!c݂�TMҫ~'�p��6�KNy,�47�X����"��$��ȄP3������]s3��P�/���^������C䱱#o�bS��<�yW���\Z2�]b�A�V���+&��I>8�߈�zh1J́E�_ .�"�2��S��*�y��{ѣ ����J�`{L��4�4<�f��y�y,2jr}�!+@rpZ��Uz���,�r$��;�G��^������2��	W?�t.�E��ƻ��G�*���Ch�QO�s#�.�M{I��Y��ZU�*�^ج�*�<@���g���q�M�K�6����DAk�;�K�BDR} ��3�?����b��4��'vo���>Q�� ,V_���\�>��J��ovͫ�  �_�1�E�[�.ct�5�{J}0�����;sB��腉f�G������E�?�!J~�6.�H@1�U'����V`��J�m����}��9�lLڒ@5���Z֐�V��ł*�N?.'�ǯ[r������Y�l/��������I���]"��������xTi���TxX��[��1x$~��O��/ O��4^�Q�+�B�8���u��[�2�����"^�.D��Wϼ�D����,9�_|���ǋ��Z�F-M�MwNI.�ު�#�X-�?wRө]/�R�S�>�-�~�=��B;�8�J������6rmi��B�*>@��۵8H�Wz�.]�Z���
<خ�d��AUo��s�Z�����&C�>����q��R�����Vǫ��B��rn�>yO�]���<s��X�&�KE�k��9׆�G8�5c�^� `3c��-�����^��]�D~}s�������̀.p�XG��^q���Uy���Ht�I�O�(�n�t8���g�א�n����-B��	�;3�x9_� �>����"��ߒ*"0���/{��>B�[ڰ,o�A�LM0d��Iz����q������b�S/�ƭ�[�U���%�Ј�ꑶ3� ���'�룬_�5"�ѥ���~�qJ0S7���,oX��	�s���-\�_��=��0���1����G�������?�