XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{����\�miaJ���rw�Y�����hR7b`	��)MiZ6Tk���Z#0�� P�!9��6A1;ځ~X���*k���/���&$��Q�D�{��*���	[H"L�A���0�^)@�nF�
)j%D��w��� ���:�W�%���D��^c}2b]6�4\�Q�����T�@�.-�`cLy�+��	ы��Ż��]}��!��O����A��<-�>�@�AV��	�q���籥l�On��c|�|�m��z~��Py�j��$���a)f��`�C���Ra��^ �	�g�7N�A-�gR�fF�O����.a �}(7�n���	!QA�El?��&yb�L.}�T0~���<{J�x3U�k=��d�t������x^u�+��>e�/��C�P��������W6��/�c��u6x�t��=�G0�K�橍R����g)���>�*Ym�d�C��O�
�\���Kĕ����H���*{���0}�o�_|X�%��لͫM��I)Wwn���f
l�e2X�`I�Z@>�=US�1���˖��+A\�/i	����V}y=�t�A�eHv�Lp�Sm��h�wb�]�`��ch���8.e�y�{j�`ܿI��Y0��ȧ��r�����V�}�qǣV��v�s��e��z�NV�Xq�q)�4__t =^	<N��x~������3�mv�މ��RFn�/�'�?}�M��ħ̞W��Jb4Z�����]�k� �h�{��d�XlxVHYEB    3b09     f80�B<���TrIg��{
��m/��:�U�E�`hک��w�ھA�j�>?P�V�_�ޮ`����)��(6�Dusɩ%n�=޹b�ֺB6f�P}��L`k"�SR�S�����S�~&�8d���s�,z��{�O�cs��ԛ5`���O[o�a&QQ[A��
[s�0�_���B�����Q1��*��*��ir�D�lۓj��l{
u�#5�����J!�걩J�"�4�۝#,"��Knh'ݚYج�<��47��U��ug�A��]Y��q;�������2������(�[Z��Z�i=�E���o�k�?J<��\?!�s��؞��5��]0[�w��nG��JygcN�|:�?u�T��tcPPRS��<�\�[��)PJK�$rE��"�zO��@I)p �Z�	�Ռ�S���%��4����{�,�sx*n�non�[P�@���ۇ���z��E��%r�Nh  �r�"04Y��j�:k��t�����~�|4"Z���̦UX�d�J�8���;����f�)Bs���i���iY;��k��HO�:)�~gE�f9���s��,ܚz�G=c����6M,:����l��Ş3���'z�[k�?������'d�I'z7��v��_�C`-�����i���{^ZHt���]�������D�Εu�+�e�������}�S�'����C~�
�/�a�ܾ��Fϝ���%Y� F�f�\P�A	���<����7�IީMJ��)`
Tkfm�3�lI�nq�9��^�ֻ�oK�rBr�%���0|�d[�P�F~���EA:��[��H��� ��bHuj:���r�����r�@� ��n�W?����RT��I;߅����&�}4��❰�)L#7D�n���v���w#���+j>g�\ro���Ճ}��r(��X�۩����6���'	6g���Kx R͓*FA����aO�2)I�|�^�/c`��s@|6�?�X��*�X���^8�]�D��mi XQ�����I��W��~��u�4u�2��a^��t�;��9�v&�~�9��^��:���s�p�/03*%o�'���o���>IRj|$]D�v��p��\/�4�qm7��C��0�e���'��� ���JfV�?�������8V���;6�3V��!�6%�Ùd���^�'sm�UJ��ݰ)��ա{z�k����#���Pq�V���Mw��y�	����L4���[�G�����[�WN}�dd��l���#N�L��H��j�5�q;M0{uA��ǒ�)X~�=�c�D��ař�<��xO�V���j^�@�f�28k��CP`l�mh�K�[F%��e����"��qx�7��X�t�A�|a��M���N� ��V�"ŕ!�y��1�FE��h�i�Hy�L_�fDk��/O�fi)�7L�a��EH,8�󳓋R�E�#�gWpH#{�n�%���ڂ5{�fG�[ˉ��@Ê�ɗ:�	m`��Y:�BծD6Ob�ȡ��ٹ�O�1�R���Ӌ�*=9�
߬Faؙk	%� #��!:=f�ݜ
�wb��aʅ�J���n�C濽U���A��:KT k�Bݰ ����]�t[K9"n`g_�_g[U��3}�﷏L-Q��N��1��ߓcUC����y�KCU�u���u�R��C^O W̋�Յ�s�y)H��Ź4�KV��4N[E8�8�~5(Uoڜb ۺ�8���K�����T%�RZ\z���0?��!TCkgrx�$ٽ�S�VSL\)hݡ�qs"��m0�:�Ng>O�S*,�27�M�RkK<J�<��h�>�uG���)�&R��Ů*C#���	�4�Ŗ��?|�P�#a�p[N��`����ے��~Ѵ����^O*D�q ��y�0*��g������f�܌�_����!���B��$lgH�RV��Ve��Z�J3����*�3��U����ڭo[`�U6��r�zd�u c��G���o�qc\!#�YǤ��ei��z�2��*{[ڰN�˲kJ �H67�����T�]����bJ��d/y�ӓ �{#瀈���]|���(�����X!�, վʜ�Ub1���n>��e�o��{��.��6��#լ�Ѭ}T�v.יc���J�|t�zRS�,
��%����po� ��S��w�ض�X|�,ʦ&���UƤ���z+�ګNO�?-��+n�����k�:H�|��V�s�Vm���_Kaf�3��%t��8���F	������á Т	=�%%dX�S!o�+`��u,[n��S�UC0����р*��&ׄ��|cH���Y�웉u����|��|�xk
/I�{���ڡ-�%[/hߵ�s���w1,#6���B�h�11�����T�Mk�q(O�}��_�K~����뎮.]��T#�%pfQ�		+BV��rs(�;n݊�Um�������(%�S�~�;�ww��l��6/�ٵ��m؊jo�U���S3!��v$U����@XM�ڲ�A���P$2�.�~Ԇj9 �uC��_�\/��Ǜ�w1�$K2I(����c�~4T��a1��r�y�"��$�Z9Wh5�Iz�|%�QFO�_�?���?��D�)�s�KHk�/�=y�7O��ʼ7<WS����T�>E������3%>��E�d�ط$n�{IO�N�7�=r�r���F�࿆-�-E_$:��Q�˝�T#PrwL82��b)jZ0,%p��¢�wm���m%�.8��v���N����R��N�L`>	��k
u���i@�����
�3��QLrv���Hڮ����P	l���Z*J"t�&1���ŘB�g�r�d����l��һ��S��$�-�LE�����]JU7�P�q4Y�P�=+���6s���UמP����1p�"��L�9�~�`���
!�bO�����o��E..��5�)i�L����c�VxW,b�zZ�{,u)q�z�CefUb�=�>.u��[=#�Ǐ��bu&AM��CZm�*;�p��S$�+a9R)�)h����uڮsJ��>�`G��Ԫ���z'���9��Iϴ�����M'��|Y�9��H��"�9�+0AiGXEBÙ]V�D�����qK��MR$/!��ժ��[u�k��,wete��� �~;n�rk�-�c��M#���e]�d��&�@��|D��"f̑��=�0���jV��|�|�T��hp'&��p�s��h��o�Щ�x�Eh7��~��~n!\�"L�Y��w��v�a*������^�*ɫ�xQT�fXlqM~%������	���fG���~2�g��'w.?0�$�����?/�g������Љ��P<��/;�ֻwi��±�^����~.�|3h��+��p���a�A^L�h����}��ot��qZ�~����]3�wR���������iSIJT�:S��ק��t`r	��ӷ��QW\p#X��I(l�֐��{�|�#�ƭ�MU�ONEx�CTk[LN�@�Y����`���А��G��N��<�{�� 7,Q�����E�Ґ�!>&�~�X��d�)�%P}���|rhw,�����/��M��O����Y�B.�7�)vOI�'�<s����2���L�~�^U��?On�������B�kB�����^G�+����+΍�>�
d�?ŭ����f� "+�8� **����QL:��@�+<�hۦ\��j�v�n�Z���vY>o���M�B�� ދ�+BI���b�xT��r��ٍ(촺�s�:V��_!ń�&ͩG��������@\����s���5���՗����r�C��O���L}282� ��y�c:AVU��B[��E����X
 �n� X�����ͥt�16��X�u��c�@�WT�C$`�]s0!q�&��	�ir�(P ���k