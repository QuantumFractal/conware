XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2)�CX�M��wHH�-�f]�w%�k�:L���+��n�+5}G�o��]����cJ�H@vڊ\�������ML��-����4���cR�K���>~���~\J۝����B���'�P�r��GԜ����?�	�s��y��h�I@��[0�i:��s��E쨛�!�5����l��D�$��k�bҒ�r^^�'2E�}���[r�ɳP����4V�[0
K��w,�jK;-��h%T�vqw��(sVW&�}"ҏ߆�|'S��9C��M
*�@����̙��A��ԑ��?�b�X��wTz�{���	�"�,�s�S(�mK/��^!c�;�y�H�>��4�M1lɄ�fe�5��۳�FN�Ŝ���yѺ�J��&z	׃u_��<�Աޮw���bٗ,�ૺk�l�c5}f�j_�I~��H�Y��S�l7�%��S��ɪ�-��n�U�Uz�j��
U�+���گ$��^�\>w����LO��poBU�r��e�mgzU��(#�z�V틡�p$a����t��C�B:p��e-�.BWjW����=3Щ}2=G[����"�q�W��{6̄{��[P��Hk��{��;��L��\�d��h�����9�L�tM��Q+5n.F�[���	��pJ��$R��oǥ9��}�]KO�9��b����E���v���n�fϚ/̡�Og�۴���O�˵#8�D�/~؛�Gsyͷ��~�s���1�����H��@��D�L��ώHh*��e8����IXlxVHYEB    a037    1fe0�?�&�Up�n��|)MU$�XӗXBL�?��J�^�_��61��B2�KTc�ׄku�rZ^u�R���C�Q��M�*i�L�� �6̅�͚��6�łD�햀-�q�f�	���Vs�2��'��}�_v'q�Z��){��M�lA��8�_@c����zaGE�O�.�C�Fh����s�
&b��ǲ\�E�/��R�X�}����
��?!�p<K�AT$��q�g&��{+�?}�0�ϲ1B�>V�=����]p�Ǟ_��z����7�Ha�&�G`���m�	D�.���q?��,#�	�n}�8b��n�ȇ���҈��e����F�}2�����3���5j���@@{���qO�LV��3���!�y�( \\�Ta���=�D�C����q�Qg�B��Z͐<9��nav��UK����\[�����2�W�CP�,.������A/X���E=hPm� eE��P��
�nUj��u�ɉ;fQ��J�$m'��S�>�� ���4��ms�H�Ѧ�9��Tƶ��U��Y9�\�X0�ʨ��]X�����
�TƚW;�ȗ�޻��3#������fI)i�GEN{U��7CL��_TN���߿>����s�n��&dҋsms�(_��T^q��iZ��[��PYRn�1��)P��{���
�(<�j5u������9�-�B������A'�V��/%mel��!��W۶�{0+b�4m��܂��A�&l��X��W^�?c�u�Tx�QU9Ve��3���
TɌ3�E�x$�j�+���U���|�qP�s5*6� �g�N6,1؏w8bi� n�����Q�N�.�8x��uq�;ZtA;��bBF���zb�]&N�\�t)����*j��o�,@��\D����I��hP����y,om����|%�~g�+JS�ǻfp�{����	D�B�x1� ~�բ"_̙��!�,c�GW�/���j-����\�C[2al�5��C�4�f}m���n�Z�q���f|�KVXj$��bʅ[V�%4G��Cu��̭����Nf� j�d{!���}f8�G�<$'}S����i��\���:�S$�b��y��o�Վ��|��R&�� ��k��Q���M]��
�ZU�?RN�tY��uI� zj�F	Frqx�����O���3���.>fj���5n0u�ù1���-�ZLۡ�9��V��>��P�+��$+(��̵�G�#�۹m����/����r��`�f�7���y��h�/hM�7}φ�@(z2 }�p$�����6̖tf�D$yt��ly����O\v�W��	��|���R[%&�<��n:Yώ��ϫ��Dh�PX|���c+}ρ�,���	�}��~�?��R=����Y�����h�� s�� ��7T���)�ZO���4���f?��c��3�����q -�Kf5�}~Ƞ�����'g.IV?�Vj�=���y�{����U(�����]rV��w�����R�nL}�X�Ҭ 7.<�O�ob��=��A��������7I�k�
� �Ac���A�cx�7�:��*�L�c���M�xem��@��1�cEc3悈�f+VK�B�M�"��7Uϋ�m�#��*d\�[��j��=��{^@PJU#���>�ۙ��=+�ܧ�Zz�W�ib��xY1���N@��O9�Z�٤aL���v~ϼ����<u�F��~?������m��rS���o�M�����B�ȼ��~ACW<B�5"S�*�|�DsW�Ӣ|�����͢�a`Ř��݂���i�k�kw> ��8�/!�=��=$��d3.�t��4��qZ����������J�����>],�Qn[1p�{󼺖8�<qځ��h�VPviJ3���뀨жuj�w�t���0��j#8��I�*�B��d��*��*���T6��F���k�r�V��!���q���~� ���e�aɨ�[��,)�� -����U�g�<;���P�W����0aD},ˬ�ш>ΘCUQE��џ��6ؗ�/E(�����풒�����y
JY�&fa�4栚`*/r�?Z���g:3LhP��E�E��+�)bU˞�+��m�q���ð)�Ov��=f��l�{[H�|$��z�oW?�(�c�"���w�3����=\�S��{�aJ��ӬEf!������'�e��E�bHU�VS�����G*D�����c��X�����2��)�V��#��&��@���������19T/Ó^o�;m�/Xk[��}`����
 �[R�U����l���Bd��#�D�+Q��wHs����I*�ŉ�$��wɅ%����{^m	bW��v$[j6�`��Z�״�K�7VFĦ��u���E]�ҡ�Y��I��P&�5f{|u6�TQ��$_"�[����f�u����XZ蛿��i?�M�$&s;iK�A��g��iO�/JToc2-���*�IU_�>�i�oZa�M�4���>[�,/gs�zW<7fI3p�Q�=�"yXV�/�vC9I�f�N�>�9��;~G/�0H1!*��^��e��G�����;=�H�5��#</{�0!�]�`.�E5���nv��j���Yi�m_#'e��|�V��.O�����g���S����/�co,��Ec���CN4��k�\bY���lVoƎ\���aC�{��if��8��Ғ�jBr/�5�wb�Ȓ-�1�t1�.��7(og���٧*����]�x�ǜ!��e���X\; �@���B���l��MO �����
H��L+
bZSx��	ҡJQfI���w.��zPĭ��}�����f�����C�1"1A�}�濚�l.��rvc�X[�]֐�+�.:���{9z5��֎�"1�b!�T����1��9=Bð���|-]��6/ti�/V��'B%��4�L3�(��?��3��p�P`�֨m�{�o~ڟ��"?�$�WN�]@x	u2� �r_���@�L�,���!�����{g�GA_��Q��Q.�(�;�"^;b�X��/y3&ܫ,r-��F_+!^lj�BM�h���N�#�qh3^OӤn�MpU��L_�,4��Ͽ4��O�esٌJ��"�h!�4	6������)�.�H�HT�c3c$m��D,-���)�s�iHq|�O,���	�a3?�H����q��X�`����GbPvB�,��`��ᑣ�2�$������t� g7��6ۘ�>+L��%�yN��ИV�N�%-�v���E��~���������)iJI�ѳ���5c5�j.���Հi�\��dz�� Ұ�q�~�
��r?6k~#��/6��N�է��TҸB˫�n�%YVxk��D�!gj�%n��j�J�g��J��vV�=E�n7��FQ��݂� e�_G�n�w��,T�f�	 ��߾ǣ|K���OO��+ؑ�tv@�����`���̱SS4�߱C.|���vA���:��g3UF���y�ve���K��(����찺ީU��1�,�E�g3U��l3C��!G�羠S��`�:�1^n��F�NF�^k�UUGm��,1+cK	-�H��pT�3�aI�� ���yk�j�ؗg����F��[���{����U;���q��֎z���݆�e*pj>��{��saw����ybpj���Q�>�_��6�Hm��Y�ĵ��꒷����������
�T�N�@e����tn2r�+}��F�X�٩��#�kU?��˺g�G�健�bb����5��>�1�� q��1S��ig��31�i��I��:��.GoHgj�S~����&�h��ub9~�<'�Դ�e:��+�v�HM�g���6Ll/�8���+�)��&��(���H\�u0v?(���L��+P�!}ďuS����g�K�ؔ���}o� !�yB�~+�aJ�*�{ e([����n�d@К��sX���]�-
FTt��^g~P���׫+d�>3��Pr�gX�b�D!�t�)���'�cKrl���|B{��@�__��H�B��#T���DK '�]������Oa��ݓB�)���N-��2.�r���a`T����rXZ��/�%Z"������@�
-�f��č}�EJϊ
�m+R7���H'}�콆���.uT��'��kۇx|IQD�GN���ϴ �͢���/!�YZ|6��c|4;~Q�&��7.�;�:E�h�4�������W	9]��S�1"�{X����^��s��k3�s�[�u�t�P�-��٨�t�j��j�%6'�SƷQj��5�Q��c4��_���XId*��Pܞ���4�I�er�����p]\�8��fC�(�=lԢk9���s�}A�=�������gL*�+83�-'u����[�U�G�&�����ȫz���z��y�/1�]��-���������Si  a��(�xY�+�>uF�÷�D��u"��d���+h���%!1�/g�(�u���ڙ�� ʛ��x<Jj��x,�KMJ�丌߂4Xo�FT���+��P�z׾�h�}�sZi}�:j��I693�.f0
�fEr�Vw����:���\\��pb|5QY�g�)Z��*��e�E��9+�ȈP�#n�a3l�����j���U�G�PFa��tͨؼ��^��
�B�􅋜a0U[t�iV�a�k�L�/f�.�����;)��P�uF@_	
���E;�Xz���X�'*o���4���Vz�"G��]�d.σ(������7�%ilG U2Q��z�į����=xk0ֳ��Q�3�~���?��چ��V(��9��n D��1_B+�o�ו���A�n�+b��K�T��I �|������R��+���XZ1���E����/�Xq��k��cp:�48��dg4�ګ(�1�m��(&��	t�Gc��ӑ���8�⡎�&8qա�uNc:gbM?NB0ez?b� �d�"l���4 �꧒J��/*�@�+��u�Z(t��Im�j5sȔ��z�x��������?˧J�&ʇ�N�6҅՝{�~(@+NqwMB]�� �IHw��/��".Ϲc���7�b[�Z�3���Y#g��&�1'p"������^�֟Ӵ��W�A�2{�����,�b������vBdp�D<���j.l����.��οH�1�R����C~[�dwJ��2Ԯk�`�>14�t�>`����¨�[1�c��-xH˻�z�ahu��qJ�S;���w;9A1M�A���m�e�*{��#��\�s"�?��究�hc��@����>��5Mz��Ϳ�3�%7Е/Zl��Lǁ!�E�Z+e�`�Я��Vo�v�ƚ�A#UV���R@f�XJٛ�|��`2�R�F��My�'b�����y Iey�r?Z4�^XӨa�Ĝ�>yeY��pO�1�`� ���u���G�
��o��v'6�2u�ksK���QNF�2M#g�uMZTY�չ�?��vӡ͔\����xOؽ�Yr�$�^��a#�3ش������@GW��,��ǣݱ�A~,��Y2 a�T�.��"�!d���������G�'n��z�5�;�1����䖞n[��YE���g�������(?'����wS����c[G�;
Ku�F$�w��C�e�A@{��:�b����:Kthv�6���%.peZ�0��D�H�^d���ѓ�D�uPnF@bmM��ٴ�.�������pB]��� �6���8���a�٩6Uһ�ߙ�?����&����H�Ͽ�X��)��@�[�v���Ė���!w�S㒝�I?bh=G1��3:���юi���7���;ۇ���yym�H/.�ϴ�줞��<i����(�Ft\�v���4hx��=�ќ���7 0�ӄI�'Yb���!�@�'[���?�5;50e�I�p�~ha.ջ���B^�G:`�B��.x�����>�)g�. 7���HTň9LM�
��S�ٷR�Rf�c���tT<6�s��I ޻I��'�eq���_� �ft_�l'�O�V?����js\
hB!����l��Kzm���tyoXA�t����g�m�}!��L�:����BeFʢ��!�oXg����A>���&
'H*ρ�/Kv����r��S��d�S�@�v*v��d�x�,�/�5h��f�z�
�ȸ�WXH,;����F��s\�4�D���#$��sțg�fu_�҅��u�Az�b�ȮA���!W��c&�_b,]��'a'��:�� �#�N謅a�Ƹ�����YyZ����dw�

v�i���[/
h���*�R�-�ؑ]%eIl�xW|��>��h�(v(��w�I�/��������/	>ܷ"�����.�DJ� ���\"�dB_�!%�8s�Ru�\D�� =Z���\�X�KOx��rp'����@߼ J\Y�*��[E�������3a��U�<�\Y>INl�W �X7|'�t$1��)�@u|�3V�l{E��c�_K)�I���"9��Yh|D����O��?�1v���ͤ���)���3�w�z��7�g��5�"��N��P���=0����3��d�"$�lIw�ru�����dS�����k�YjA�[�-:v��+�9��ߎ;H!h8�u��l*�#�d8�v��lǪj��N,�[�[�R(ٳ����n�=O�'_	�u]���p��0]	4� `m��"�l�Q����IO-����J����<	m�ub���H�z�q:�F�{���%��l��W�nl��X-���L�bЅe-�6��|>آ�F�2v�[8���l��T_G�q"!X�������.e�y��G|%T��jŸ�S5^ꐠ �����x �4��3;l��x8o�1�/"e�%��`.�7�⣘�--��`W��4}?G���w��|-7l���fmH���E��? ����}Բ��RcǀxI����A��ӑe�P�(���N�f�����k�h����zEp)����,���d������j��Su�ظ���]��W�V�������K��j�R�o�Y��x�*Y�����+�Abb6�r��]ֱ1^[��}`F��������4������V�l(����Η��y�ʡ����֒B�6��M�3|�����I���;bv������[Ǟ!�t��_ڏ�(�P �);�1q���T�;�,Sx�׾���T�+6K,�y��D)�㍈�<��P���S�BS�)���Mm���hqQ4vX����Px�d�̄��iîݍ���*��i��4K[԰% ��who"	TjT3��m"I��e�u�;#a
[���7;j;;S�6��%��/i� ���)V&T���޷'��'�A.�������s�e�ľ&�}�7 �����0㍖��XwW���3�,˛�7�]���hKo���FʐzF3��;Y�0�j!e�,�T6S/�e�R^����so)��aqS{�e8BQ���N~v
��$i	�����ө?$>��jJ�Q�8��e�y]�Gj~�W@[o:�*k�vU<�_ lYU!ݴI�Q:����,�X��z�������O*�`��ܫ)3qҬ3s2x�߸]�+}��7���KD�D��+�U�`N�y��K�Wе���]�~|M�'�����X�ֆeԐ�'�S��A2���%{��W�������*���lȒ�'?0D6��~L.���:�jA��]�+��܂/���n99�̞��-����DA������d�+z.���4FJZ�ˬ���n ��H����>�h�/[�~zȃS��Ũ(��TЯ])�I�뵦�)���� ��b)�|�w�Rdkɔ�D3��P���0IsrgS\N�M3�A�m���a��&�5��{�����\B�-N#���E+�Zl�R4��Ā��.9�n8�n�e`�C������q�W� �h�t3�Al<�[9R�Mn_�\Q36s�ݥ�T��6��:wssヌ��LǢڎ�Ŵ��)=���I�7�eŎ�|�Y�%��{������D%�,b�K�E��2�"G�JKQ�,f2O��ey��Nu�B'����