XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������󈸐M���U��t�ŭ�� �^��3��r���5�K�o��-@.3�߲�{�zZ/R�1 �3K��?���D�,]�Zn�=Ȃ����v�^��7��~P�)�2=�S:0���U'�,�$V�T���`�����r��3�a5#z��͡�g-G���+N��-�u��ץ�wʟ���y[o	�\����HE��Gi�a��ݪ�{U.4ѯ��ŝۅ��m�|�3���Η��C�3��G,�4��Q$��Q��bkW���c⋬.�u}�;�x��b}�B�'����#�ݗ�%��uJӒ���	G/�$�)��x���Ғv�ɾ��6T0�]�����e�}�&�d��Jܵ�Ah���f
D�>˙��v?�Ǒ[]�b�o3J��]��nՙ��.9]>�G��o�U���W~����D��%}dˈR�<rW
���KN(|Ȕڷ�qw?�^��VV�D2F�}���� �w��K��<g�ŅԛI�7���^�K\G��9��� ����N����G�3���-G���7��wkB{mu(��km�
������5�R �l�"k���Y���ʩ�!��A�[�ٻ��V�b@�z,-�����uR�o��"7�V��<�_Qlß�O�/�PW;JP�fu�,�(@�+��Y��kw1�.D�}���n|6�'��1h�����d �w)+G0}���'CW�Z��ɾ $�6TD�ٜ�������3�'2V�I�2TXlxVHYEB    6014    1840�1���ztV^��X��aߑ�?�}�E���ѕ��gǈT�����Z~��R$~��M�s�2� [W��`]I:�XW�:�K��ڊZ ���t]���%D�%��ƀ�N����F��j�N����f2�� K-�uG]��R-c}gLV�-��F���;�xc#����������z��v����Q�w7d�5I��U��J�o����nlˈ�D�������j�B�@�h�T�e���T�&P����bD1� ��f���-��j�/��M����P]�sq{b�om�Ћ_ϵ&�]pu�O\�U������Ξ�Lw��3��׬S,����C���~g����� w��*[)�7����,�~\\!��`�ƞu?�R�w�9ק���U`�Y�FГ��\��Ȗ�-C�9�]ű�հ=���S�yͺ`�|�o
�������{����ъ�A����ճ.m�Uv�oo@�k�U�t���F
�>�MG%�p���Y���T�=Kjb�V�Ao6�3����D��.�i$*� v�UF�KN5�N���^�:N�7�\�O�H)�+�ht��~ Fʩ:�.�����	������T�Y��fҲ����9�������1��:���P�ܯX��|zǿ��TF#_�I��p;0bv�j���fo-���d��E�EP�C�����N�����8p����/�i �-�]����	G	�,=��R��������Q}7!k�m�i�h:���iB���
W��y�md�T�"qDN���6|��h,�/��Ė� ��u�-˩w��@.��L�����ݥK9M$~Te��bуsXyȞz�p����J*�Ύ�����<��%&PmG{���/&���mK�8�8�|!�}�hW�L}`���%��7K�#-t�?C�	&}+xf���3B,��ޟ�p)`e�Q?,sB�[_9��^x�X���n|���۲��Z�#���M�P�,���v��+9���,in!�E��V��+�/��E�,��r M�(���g�v�'� �&Ԉp�rԊ{��������(e���vf2�i�RN�W�=k��H��Tq�*�f����'��8Q�9ў�8���C֗D�/w�ʀ�c|Ud[~��x��FlRp��Ɛ�}Q��s��w#Lc�(+�^��:r��#P܍���#�l�b6��0�L'ҩ_R�89��]�s��! �[?k�NB��g85?U����`����96P�QX�ݸ���ހ?�<�w�Du�T	���v�0���~x���V{r�=&�&WM�(5�:Wj'GȚ��|�%^�H"+��<�%-��9ɪ?P`�+�}��s�^�ӯuA�]����"�5�JI��@���K�T΁�i���$Oa�s��s,|��V�Xl
Q�G1�x��Sd�̏xۍ �2����󃥩�$~��_�C�Py!^:�����/Y�ډOW�,�J �ewX�3M,�rAJ��jϼ>럫^�t:a��G�F�Z��h6(�ov�w���B�ХyP*� ��?8��U";DA~�$<G�ip5�`�)���7U�g ��H\���1^a *�U%�"�D+&Pa�!Qm���W)�3L��ѷ=g0 Y��-Ĳ�f��PΟ^����H@�|q�7�����y�����Y��|��ʺۻ�dc,�.6��f�Ā�Ḥ�Wo���Vp�/�w��`�I��$_�(&�lFy/���G��_6����G<�?e%�l
�ġ���0�b�!C�j�(vp`�V�x��$g�Gv4�G��y��-臯(HV�]�e6/F�	��\���<-���_������z�QHwů(�<�U#8>O���ٮd�3���`��1�5�$�u�+���?����+�L2!Y��}��\�fY �\���O�9����*%�}}����/�A>�$��UΊ�O0Sxl`mj�u��<KY[<Hd�K'@U�!)X@�NDK��.��V��,�PD/�PSǓ�D�VFJԂ�yDǘ�&�ܐ�s@V�,�P7W`Go}��z te��\��1|�(e���rKnl@��!�pj�tzԩ�&�4FNr�0ĥ��]L����;��3(s�7v��0"��S�@�T��K� �	*�ِ6N6�r,(U /�'�{6�t	��_-��,g�[�W�y�'�߳��Ĭ�H��9ɚ����ح��5��)����3�p�ز�$����5e[�t���մ��I�h���)�������hł��b�ӗTĤ,>��Ȍ�hFU��rpG�nH/� R^�ηʢHFqRyx�M|"e�xv>J��Ԏy:nVQ7���r����.�
NT�o�������> kH���W��5�@Fd����x:$�0Quڔ7�K���i>���]��C�z���ٰ5\a�,	pd��O/T�G��TB�0JÎA^����������J��=���Nr3J|6�ɭ�9~�dZ�)?t"KJ���e�h�B��/�}�SI<��T�e���H�%7-o�k��4�p<��bcd㻖�K��N��(<N�a�v֝$����^�F�2��=6U��m�����ȥ܌���mX�%/�:��}Q��6x��a��0N�h;���NrS-C[��6ӥ<±���׎p3����ߨ�%*"9���E`�K;�؇��8��w��+̆m|�#����J�ma���Dxǥ��%zSe���'8_!>�J���z�C=s_�����<��/�L�;�x7�:��g32��%����2���(�E@N�,�c"����j����\���B"7��݆#0� ��]G��O�����^�.+��$��j�6���Q�7u��-����
��%�/37 ������ �=Ep"s|4��C���D��A�����S�h/�S�]A���$��ȹۂW8���u1�=)�#�a8�gk:	�ȤTI��ޭ]�f��XPw2����y�B�w��FD�4b�9�\��:݄�O�
"�y�����X���auڦ�<U*~��'y�L��io�TI�d����a2u�)/�H�ף���n�a�|��^�Lٳ*�)-}'NH���x}(��$�������C��2�����$�7?.2`ƹ�F�|���R�崽:�w���'&N|�s��6���k=��l����(����.E���TMh�&����;��zXp���+����y�J��D=��4���]���}��B��n��/}C������n_(z:;�&�3��9�d�ۍ&�?6֠jx��P�u�װ���n{P�[�VI[1�]�ԕ�Qo�7!j&<�n��N�+�-��x��,%l�K��g�e#=���U;!+E�W�nܡ:䗼�܂$��_����А�b��zșUE���㣵r{�4c �"����Bz�AQ�HnF� ��r%��lV4��k�	* ��>p�ax��Wy��>�;�m"O�>f�f�qu�����&�6Ɨ�scK�o��	3u��}	�<�:!��v��K���L4#F(3�<������|�7���iw�������a�ʨIo���-�<��zPr!!?MՄ>g����߆Gp�֣L'��+'+�o�_L:Ǯ9\W�۪tz�'�N������a��Uå�����_V�>l �����Pa�_U�Y^������Q�����Ɉ3�;޼�#`��Lq��#��mS'|���yh��0<��ޜ���=�����W��v6cj�^�M�����������S���� 1��*{���R��)���PF��yO?}"E;Z�#�����0#�l2�&t�g���7.lo�*\�x��I�oj�� BQ$@���c�{zVO����`_��i>��1��v�l,���sV8�Ģ�u�]��	��#ƣ�w�N��(T�H~3[m	�7[�JG�ʋ�:L�W9ę?��W��>��q���7�S�ND��ȩx�����c��ړA�a�cM��@�Ă�L��*��3(m�C����W�����4kJ~N��Χ�4�Vٻ�Pf���c�����)+ib�!���d˔��|�}�My;a�1G�耔�ͥ���>\�j�J�/�0HƑ%������a����3���
b���Yl4Dy�L��nG/;]晖c/1�0���a�y�����$� 5��t�R ��eIZ�����:�M�GSI����L�x��%+ߐ4��`T��9ޅ<�[a��E��	�"�8���LR�5r����u�u�i�HY���-���k\e)�v^r���Wy8��}~6\��^T))36�7��m0>;Q?�~b����y��-_8<���s�
-֞X�}o*q� �cJ/#��}sG)����g*{��۹֝�-y������g���nG1(�_���@�v7Zm��C��U��0e�pB�[#�D����ҩOf��ur�]3l�s������{��Y:̺Y-=����>)�x�L�S#�X����sޟ].�\mi1@ޗ�ec������ʅ�Nl�h�^�q�p<���I|"������7��k���}�A�!Y��~�mV2S��3�]�0�1�@4gU9k~]aϣ	���\c����/*��~�.M����8��s n�Fw�Xv�(����O`+�rk��[�]��Y_���ֱj/��3\[t�Ǎ!â�%n�:5=Y�ia����8֜��W&�~@ժnKN�i��,eKl8��X���M���p2�N�|ņ%��h���ie�S�~�hٔ�N����z�ZҾ�M�.��> �^n֖��g�.������Rf��a> g|�����M��T�M���N�c$��щ�Ζ==�k�t ƭY��*7I_AqO�.K\�?K�%b~>�]�(�z�8�ɍ���j�-�&��U�&b��,�Δ�O ?�����;w����k�)*�]�(kѶ�a!H����NKOԟ2%�u��Y�綳�\N�J��?��#`N��	�?��g3Z��L���T�����?��A�s���^$���}���a��/����2.XYh�	?�a����=�2�v�]�)�.!Xy������3"�m�"7��2K��O9��G?��xǇ���)��'�B�h���QNK������E뇖�򾺹ɣoNB��$��؛���G�1�$_~J��K�Vȭ���r}�ƘW�k�8t�:��V�`%�K�Z�����S��w5@{��X��w��!��B>�.��Խ��x���������w�=�5�CH�"bm�80��SS����9�bo1pI<���0뱣rR��'ǛϬ܎߬'ƞ���p;.��ہ7+E�U S`01|�
���k�a9�)���Ѯ���q�Z!����WBg�F�C��$��|���4����M@��\��Hq�DPP%��!浄x.�6�
$�_��:�����V�2]^���XG�7nܨ�3,CDFٛ��W{yY;lxF��%���H���
˳�~�I[�M���m$�|��8j��q+���Ψ[���𣈋#��m��Tb`��Z�C���W�ܚ#�����bM`��Y(�9�	�nC�'��()����Χ,�(aH8�
�sq�W���-�ļ��)�<�|�������f��nw��E�F�&�/!�I�E�EZ���C�O�ȣ��f���D�����!��"z�&hu���1�nf^�5V��Ic0M����a�j��0f�v3

�߂��%�� �Q3�NE���<pq[���IAB�N�)�b�I;�4�]�8��15��D�@���2��v���7���`��.�uc@ǿM�=� ~`���r��9���_��	�i���-���5ʉo������a"�!. �n���V: �����CZ؟�J6�
nַ ���Z@��]��Ƙ�=G�]�Lx�1k�.���B����Y�y8~�&�C�a �R,��p�W�b5�C:%P�ۚ�;)<7%�~Q�:��\�<��Lg����@c)M�l�ڄ*[�׎���p���?|�w�>b�8H�H�B�u>�!3UW��o\��vX:��5��|(4����ہ�Q�ڮrn>T7N �̶��(��O�OaWȥ{ӎ��?݊#�ֈ�k��I;�aW�X7]���-%���@s>�[qn�l*n���H��=Ú��M1tl�k���8�