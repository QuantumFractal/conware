XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���xGe�A�O�8�8YI���dl8@j�x{R8�\l��Z?�1oO�pk F��C�)�����>B q��t�uȺ�=r�1Z�� �U�.G5sZI/)��=	H�_�8���ӛ%�g�bd�9;>)~P������å��96��X��}�a��.����`��2w{�ը�(�S�Hg�cn����Ӆ)S͙QS����@m��T�qN@)Ɂn�#�q�b��%���-Y���R$u���Ԏ㾆�>w��\Q��-�x�(7n�oN�����w�;�_vU�l�3�LpPD'#@�8��ܵ���T�(r�Ӂ�2K�Q�څ�kc���x�@�$��1����N�K=X��xWdM��?�Q�5Y&�����3�8T �y�t9}�;�� �TQc���d�nۈC����, �q{Ȑ�NR�d�?P�q5e�MRʎ+�,�3�<��l@N�XK��hp5r� թ�rEr@�χA�p�m�s�L������D��k��	�5�&���lG-O�2Y��G|!��IC�.M;�|����IBhN�@�k3����
/ߙ��C�N�J�;H+GCx�p+�3�;F�µ����W���^I^���8������|�=�z]W!��VoE� �IS�t���6�{��و��x��R��-�+P�?T��W�Y)�T�ϻ�$. v"��d�R�V3"�<�6N-|���p7�	I��W4���/�p����>8�߿#�Ԉ/XN��i�
�$1�ּ����H&6<�*sױo�k�y*�z%gFXlxVHYEB    6346    1790�����"�`Mn1�)�4z�s�8g|�Դ�XTz�����`v�xE�{��R�(�ii�w�9f�D��]2��V�<_\\�p֏��q� ��{!G�.t@���V����=���1H�e!>l#�_"��P�B�w4�`�i���r�tZi�aaٹE���IR-�� Y�nf�ǈ0?&kks���h��uѡ�B����?��L�����c�Ab��w��m���:J9���*,ŋ~ꎛ��Ӓ� 3�l�&�_H�s	U}�?�|6?؈l=ƙ�Sy����vj�m���u�ƴNU��U\ݥ�7qaC#{���,�UĽ|9���m`�@��u�:Z�	��(G�J���7l4����N<����Je0H� ?�a6���H�Yc(�.#�@�f�����2К����[b�鲁R�W1�MGd ����8��v{*]@��?p����?�N�Zb�OE�Ѵ�������!΃H�?7�05�=7�Y��4� �#s乄�� ��wj�/c�;S��y#{A�u{�}�1=B�@�Ol@U0T�O+�F�gռ���R�6�;�_/�����hL�/�ʨ�J����{�L�%�Rd'�U�L��4�>�4R�or��~���׌8��1��xA��� D��a洩BZ-c��22vd�k~�*Jt�@��j�TZ:9=p3h}Ia�l�
�0G��x�
���d��j�����%��o�Pʯ�PtM�P�y�w�3m�!l�h#lORXJ^#�E� m�d)3�� ���+`5� '*�M>�*���(��~�sZ��d:u���O��îR�x�<Z��ý�T�-�/�jRI�s����Y���r��'�|�J���<�k��
D�/�}g(~.�J���3��i&��?�8&�*����2_W�~���ǫ�^ŭ� ��k�{�}+�q8ax9�Bg�-U��=L�*�����};�D����
&{�Q
lUZoI{L�5-�����.�ް�6���1ȏ��7����k�U��6����v�恉���e�~#���]���Av�^P�����ع�	��4C�Թ��G�{K;���[�T���G[|S�X�F'xX��м�=G�����P�B}�=j��Hԛ2#.�7�)����A>�	���,W������$�B� ݔ�c �òT�����V�o�6�O6Ì��t�J�(C��ʢߺ��,$��� �_�iF�g��m��3��o*�7+��T�z���A�=�9��嬈��Id���6�¦��q1��=�2m0y�=DB�+O�s��V	�dK�ky�#�{�kɥ6K�ꆣ��ܽ�@�`=y������8	{˜qF����-��]��N�O�+���Y��d���m�cW�smS�Ҏ���ۏ
*�N��o�����5�.6-�L�{��|lS�]��b?���/{c�M-k���U��y��&�兔�4R!qbǮ�Nj�9��e�xnP�U|6R@��X���8��
�t�qDC}����8�sJ�Dy�&�cL������wE��������m*@�z�y_G�>s�;�MN���1���� �:��OJ"��s����E�4��oK�6��h=9
�诉��2���?�����a���O�)�E��o��c�"�g
Z/��[�5E�Y	��6
���5�'�atu {,~��.�ۚ��������7�� \[պ��3b�� �,�Ψ��c�5�#kFG��J i^Q�f)Y"��!OR�/�'a�Z�w3�	�K�p�I-��uݶ,J"��H���O��C@ݰ�QWi���Ε�1��ߞn��C��Ӊ8���@�a�>�l�!Jߔ��k5}�~6>%Z�by�勖|8Gt\u�mq{_��l���D�[�U��n�|�����ܼ�ޱ����F�o�ө��vQ�n�!��������s�4�*��@�?p`��v���{@�K[s
Fm@`���=�iG��OV�B7�,U�u��4�\�w$�6$i�$��l�'u2�pF&��EL��C��1{��I�%ȗ/D]���~8�<t��?J�j�U'e�~X^�����L�*�ߜ�Z:����(�J+�#S�Q�v��zaްgUT�FM}(,��X�<;O��My�T�p6�����^���<����9Aoc���(�#�0*��Jᩆ���3����S���&��[�������L���l�N����B��"���lғ�¤d�9ɪ%��sPĥ�0%f�5� 1f��tｄ=������"�����v�u��O��eĦ��8`Ǖ`�6"g�s-U�bk��c��F���O�o@�}FD�j`Ŝ�z�!���o�l��*�|��0|;��:��[�r�/����pތ�
��[f�s�pG�ȸp����b�r^����Qi(�a�ȌQ����;jx�̨�t�d�"�ͱF� ���x��a�e(O��A��3���hY�|[pQ�*�s9^QR� �P�Y�3mݲb�4M�g.��ꊊN*���/�!.jb�I<������i.��g�< ���[�I2���y� E&Uٵ���<FJ:tIp+���:]�X]U�F
L�	H�"-6��U�BC"N�&8�nyS����)�m��Dиt��$L���A1ߧ3� E_�wR�;�7�-���H�%96bWU;��!e�kL�������י�+K����A,�����c �	N�ۮ	<3A����BF�yv+Y!X�a��.q�-iK�+ɜ�Xt7�H�~q�ł��0]���dx�Gj#Ȩ�*''���fdD��_���~�!1{>�mʲ���tY\3��=��	��qVw"�w�QpX�������@|�F.~1�K<���&�4��/j�Bs[�3<C�b��MLr�����MU C�v�9r�̀I.���߰>�,���G� �$}*"� ˒����,:B)�O��}\�(��k|."�
�sܼ�~�mɉ@�=�o��r:��p���߶��>j��t��Tr��Jk¿�T�d��zA	>1�4/����"�����b�g�B=ݥӘ�gƷ��ҐvL[���{1�Ll�YH��@�G��e�c�_e�J���*u���@y��@Ƶ��	�+%ӹ� M��8���R���WW/辚0��H	O�Z����l�A��i�����ew]F�c"
�1q1��F��S�Vp���r�J&�5˧a8̏;bq"�=��U��/$^�_&E� \PdB��@[�J��ͽpۼ�@
��jɣ�?+9N:S(���p!ON�O�(�*L�T��0�j��A�q=�j�b��M1�E���򾶝z73�4k����$���q��i�e'�Ir�M�{8�~r�P9�EN��JA�@Qt���H)�`^�	�����_(�|)�CD�K�bFy�/e;���y��U�����YX�����TXjv�q�%9�Znl�&��e�"s2����K��cȼ���ځ����jƘ\<KӜ�[�ߘ�,���"���N����֝�$&�u����$E��z+��̬���Io<���_jV�К�P��'����q�H�#W����N��bB�ݡe�Oo_�R�ϛ𚤤={܁\3v���Z0�XJB�(�`�hh��?7@���_���.m��M➲���4̬�[��1�����!Ev����z[SQ�'=��\�Y1�����t��D����42�~mk̨����U4~�W��k�����Ӆ��z�F�R�͟��B#\I��X��?�N	C�� �%�8VI ��W^T	*�T`����G���[��N�R_}�\��d� ���ӫ��wP�<������[�fRr���k>�D7mY�^��pw��	W.����͵��k[��y�8������鈨������#{�;�G��0\#��Ӧ��������&�	�K�m��K��I5%^O���I��+��҈��mz�䊶�V�x��S)�ε1�O���I7��>Q1��{��K2^�7xE�iF�y�w�ٯfP>òu�
�O!^�ڑ*�wy� �ā�'����֒y�\*��L�l5�H�-r�����:���|��a�������睉7�1��++_	cto���HnO�ۆ�(�5N(˄Q"�	�,���Y>�*\�CYs��;����}[�!�ͨ��/�<ɽ �[%����?6ֿ@�_��%�ʶ��q)�k	��(h��dA�#8��Pvf�t�qL��p�&��E/���=�}JJ�A+��������Jx�Rp,�p�'��7��{�3��0 ����d;tޯ;n���O�K����"ћ�d�F;[@ �r>a8>t�� }⭤��
�仱VC)F�} ¸�*O����V�F �e���-�u�������*�>���i��Ԭ2J�]GF�$j���
�2`���E��r94^[�B~��G2xT�e`�����Y�
�\���F��kTޱ^"I�P�~BZ�-��߻�&�1}���~�\4��~��b���p�W��5��X��$�Ec�Q@��������ځ1�:�Y�5`��� ��ӱ�V_Jg`j���sv��v�$�]��z�7KQ�9k�$�~��:�W<�$�o�`�Z���H��5�t��J�%xeP@�rso�QB�!��ָ��Y^��;o/'�q|شn��A��b�L'U�.$:��͏� ��j5Z�ѝ��¼\'����:'�4Ik�Q�9�����`JF}����_����K��pH�<�-:u���������+D�:�$���p��xky���ԗ��2�|0R�3f���dP:�O��I���
�$Lu�Kz@�r��1/Ӵ��z<��!u:��X:����+	3�9<�kh���d�cU'���~�Dwvj����{���X�H�/脃�	��4 d2�,�9��T���pb]�d�b���x��x�� `���l��2�c��{���jZ�T�h��#͸����`�[����	�X�=;+���B� ?����~�cD/���GM( ���
yc���6�Q��=��vQ����y'��y_�ye�\<[�.�.�:�4�w� ��u����Z�=g	K���e�����gsO�rg�a"j�z5�ܺ����\�n�����f�4��Ky�F��Wv�$�)���1E�l{��M��-�o��Y�|�"�������?��6�a��� \����������`�ܾж�jP�}
�R���Z@�}����^�P�+��3еi�~�of�G����T�Մ��k�W� �s���.}h�1M�Wύ'�X W%+ez����>����zʜ�db$Ƿ�u�m�B>v�k�#����x ����Ԏp�v�d��[I�A�3k���9#R�]�`�7��p�V�Bb���&������iQ,�?��UݭOP�zCV��ń޳�r��<G_EB^n/�#���i���i�g�]}C�S�"���<m(uD
4�.ܧ� �2j�}�C,4(�,Ĩ:<(�;���9���#}[2��<Yp��Z�����-�r��Ϗb�74HA�6�~
��1�;�;s^��gA���l$�����"��F:���V㹥���L�~��#EF�H��%Ȉ�9�Tdg"��I�EpR�ƃQ6����[�lD`�j x?\G��齌׏��cL�Y]V�����h�9���ZA�_�2*�
2xR�l�0�.��d���f�҇Ul�48�[��)T�B���$CtJ����-3�va�ץ[&C"�5� �q3B�X�@g�E�]2�r* H�v���񍓒�;����Ϧ�n�*�.sw|��#��Es�+X�a�'�t�;����Uo� �T?x�!�2<Z.���VB�,�����������{_�J�߂ml�o��>eX&�z�>��$��!���lvN���̿�N�u����D��o_��N�{��a���C���E�̿�_|�
�SZ��:��4D�E
�÷��4�p�g��h�f5��}�Ԅq�@&�U
���+�Mʿ��;r����or�����wU�T� ��8��J