XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���$������(�ª��Aq�w��Y�u�g�@��je`&]��f`[R�S,9M->��Y�e/-�2�jK�+�r� ��a ���6����έ%�X�w�&�D���)�,��(�$2��\O�z!���н}�`�ȡ�4����j���&�Θ9�B�<Ҳ$n[�f~<��U97!��^Y��M$|�fPƚ�����u��[d{��
�;�j����V�Ӌ>��
��_�6��Gγg��}�
%����\�g����Khl���@)�������] -a��Bg���t��'�34&և6��S]������$�-(�ǋ ��C�ÍǙҢ��3�~�S�U�, ��\��x���_O�D�Z	I�x�MGf��u
'{q��	K�\���W��=pϣ�a)[����
7��G>o���at�r�6�O5�3�>]ޢ�M�j}�\5�����1�Z:m�6yT)�t?t�L�˷u��Bo�p�dš-_��El������!����ix����tσ8UA�>�R�aˬ�' c-MPS�i��"�*��!p%�	 @�!����!��������Zί��f)�c��Z����3�M�I����^];kG��sezy�% GkD��iEۿD�C�]Q�5Y�hq����ˈy�QHgv?�B2�E�Cg�Ed`I��ҷ�2Z˃�|X��}�Vr�F;��<V��۰S�t�J�(�1lҡd�������Z�P8�\�� �!G֏��RY��a���a�3&����� x�žls�XlxVHYEB    3fdc    1160��ͽ��f���sA9MU�%F�z��)��R�ll�}^h�X~�����Dޟ֕�����~b���2�ݵ
�q�m����^��P#If^��G�5�M�`�s����M����;��}��P��� �0�}n�ꫵd�n��F�^*�^�M�/[�Sn��B�-��ޡ�����OiS}r����)ӱ,@�$�zCŏ�w��#�E�d����֑х�&^�DK�9��R:�vQN3˄�(��6��n��HF���x�`�BP�I���(~A���^�Q����U#�V-��9ޫ�b���"��xЍ��E��o���j��X�LM��)odyc�S,���f��#� ��Fdl��մ�<�n{Q��ǢJ�H�L*��t>��\ɮ+�I����L���j����eE�V���,��2����Dc��������g�[��r���$]�{jl��ʱق���HV��2̍�����.���%0/'�*��fS棵�o��9��{{P�W�w�`�v񝟋���WSy���Q��b�<�,d�਄�6az�IBS�r��g��+y������c��&�Ҹ�����=���`������=��c�
�#n_8hS�e�m7��9��:2z-����Ex7������6U��~AZ�)�+��jE�o��ϸ{f����Et�,W�R��<K�u�e~o˚�)�RH�0`d/)v���:�����ER	B�F�W:m(��u���k�;�6���'G��d�J�L�����sC�2l�_�ݭ�t=�P��v�P�"��-W�/+f�ß)K�Z�oa(�!��,�T{�uT�a���n��9N��/Q�b����H�����[����[�V_]� ���1�A��[�-�����A�Z,*���f�d�S��P�ϕ�L�5��_-��î�&�,�{���O�����q�mncR�r����=��+J��Z����#!�5b}��iH#X��.<�J	6�0sv�ll�����X�E���$Dg}�Ӳ}J��RU��+�?���x�Ui:�8��_I\�R�3���Rdp�b(�<� tt��Zm8�e��� ίL˿���|טi*)��i��V��p���8;;�sm�@���Z��A���N�Z2����.U��ȀBz��(`���wM�N���=^�ī�p���>��[b����+і�nt��<�h���Ӽtß�_����I� �8uF`!D#;d�]�������L�c1��AH�y�K#��yž�����KК��p
��M�䜂�_}�m �ڸ#���'��3��]ב�O�:S[?����Ip^O�6�l	�١�&r�������y��%UJޏ��t��6ۗYTR ����/��FwC��AEZ��}��s˯�\Lhj,Y�p!t5?lؙ�:�ꜩ�P���\��j������K�7ʀ�)1���9��g���w��j�p\D6~ΰ@ȡ}	� ~��|ڬp\݀��B�暴}X9n@���+E
���B 8�<���ǖ��(T�\�b �bB���o#kSUM#	+s�&�#Vx���<����51D�(ޯZ@_�W��'}7�RЛ}m�i��l_{~X��X�;@,���7���\
�,�8"8�q�)y��\E��:�6�0��9w���-l~�-��D5��0�3������on�
��JXU���7<�χܱ\69�c*E�W[��-��:[t6��n戉��Y`P�Υ	�0��s�����o��+WJO-C��έA�5�M����خ@#���O�t�iH&�#w,�v�0���i��kz��Y�M��"&���5��뉀�Gc�Kfg�*�hX�!�5�	R�r^�Ѡ�iV�d�]E��t�ߊ�iK��u\���>,.OE�?dQ � �>(�Th�$i(�f�����%��BX�<��2o�)��H�-�0��yQj 8�2�� �{1D^=Z1���T`^���0�7�����q~��^����I�Os�z]�i6�uT�!��?���Gn��&�����~���!�Kz�`aU� 94��UzV�+]|��S8D�Wsپ�̐���0Q^\`��K9��N_�	��E.[�������|�u%2ϸzIR$q���o�� ��Am�
��)}p[���P2�]؆^r�B�;���#�)t���p3�ħ �Q3�2s�����.ml������p>�[����zT�ڴ`�.y�m/�)p�+�)��D�ɭjKe�a::-�a�ψV@�/w�W�Q炟���Ёl���r?(��3��ᴖE+��gPqE�׾t��Lx�u^��z}�������V�=�;#���zo�B�2�v�))n��#��u�/��jQY��Q���4�g��Kܾj�9�Vl�KX��eɣt�%�۴�T{y�~m���W���zp�@R8�{*��T}����<��R�^�@���S�5K,H�8򎧪��drbq����U��%���w[ھ�ܗ������6��QW���l\u�� eTL3�� y�r�[:��!�(���u�mN(��O���E�e$�J�z����	#�e��<�Xp�E�	H��E��1��bp�ݙ8 �'c�f|񍭉JbL �G����H=���K,�N�K�� C�&T.P��cn]�l�Hb��ߗ�i���0:ǜ�QR���iCG�!�������D0I�ȕtI0�/����Pf�E����|�Uvc�YT�Ⱦc�3a�źzۀ_�_�m��(�`LY����Ĥէ�>����H
+�ܡ�$�=�YZ*9�^��6�=�xW"3H�>1Q���N`�~����զ�b[�|��B5F��}�����y�����������r!ެh�T��j��,[���E%��%� �/ܤt��<�鶫���pV�[��� ��_�\5E�O��P�mz�^��cZm���<�}GH����ߣoV"�%���k�G^����۱Ù�}�p�z���b��{c���q�8� ��k&�Q-�N�6U(5�WϚ��{5��b�fIS&,�bµ3�S+��&2��kSp���w,�J�"ޅ���sok�pS?��F���o!�.1��鼚�[��D"$,rh����~�D���>���J	��W&26?	 �u3���D���.X�ș�:�xt�$���83X��Ŷ5Yx=���7�׾�3�l9x��9�kQ%�Id����q��J�e"[N��N�� U� ������c��g��M���%z��I6Ϳ�ψF|�o��jh@6��ݧs\����,]�V�C�`�[$���6��G��V��y}��Nm-uvLI���E� �ja���S�ck޾Sڲ٧��ݳ���kW5������ڠ�'��W�����X�k���Сْtt/���_J�I1|j9 P�{�a����7���-�Ƿ��)}�_���[ֽ�Q�.�FG�%4Q��Ss�������W��x��U.��j��<��ܿ:��kIn�/]%��� Qc躓��Of7+��Θ��rv�n�Hw?�S҅}�$��Þ�5'����
 򉕍XD���1%��F 3LM�^G���,D����K�<�|����zGoO�F~&d�cf�R�o%����u$;e� �Ϸ0XT�'M��!`J� 
A�D��0BF��D(M�E�~�c�A� P/�e������v9��޳��3�V���� �V���mY�y���8f�"w�v^uvXw�QЌ���=}�d�@��/麰 ~�����l��ݒ�l�Qu�?�����v�yz����Ih�V�� ��Ę*ʭ���6�v�H�g�^���ɰ��Z"@�Q�k{��Cjp=�.+$���V�W�;�j�1��^9�uA"q?4������MО^��O*9Z�Z���1_�C�I��z��n�V����S%�*�s@4�vA��7J��H>�J�Ҵc����b��8E��7��lh�\h�Rp��1�ɢ�M�3���up�<����]�v����m�����9g����Z�+����;[���yZ3ԯ��^�\0�G{�q��Q�.;��B�;y>X6;�F&i�8��fTU;�Q¢p��8�d#=ˀ������@qFe��v��l6���z��<��;!#��2Ey6���]3��F�K�M�c%�������Z��Ŏ9v��>����6
��]�2�L�o����J��.��[�)�B�� ��\	��H��^�E�B�f�i��
'��
vy.��� �A�܃}vHN�
����4��q�	}�[�
VBb��c@Ǝ�&ޙ��g�N�87ʠ)�r�+�G3t^��.��a��n���5�Ic��O�NE�t�������[Y�	H'`�,YÍ!x�.��>���@���$Jb}15s�2Z)�¯d��}`�%�`u�"0J���9�S���uJ��