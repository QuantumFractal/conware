XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������`�Ui�rvՋ*��iT/�e#��'5�z�Ȝ�y1�Z���D$׵�h6֮���ti�hY�-�
H��\Pyb�]��*R�邩�=�0�C SpR�H���5�4�MJ�]�w�Yo`wo֢*Rv��nV������;Z6-%�)��$�F��锨�4�Q�mo�ř�����J��;��G����Q���hW꺗V�q������Rӡ��l�����TaCz�t9�u(����\�j��%(�I�:�rx.�C>LyT�(M_�p
��`�o;�[r}ȚV�<��@��7/>\5KCҘ�b[��r�n������֓�.��u�d\鏻}8#�%پ|Ki�<�ԫu=>�~�ͱFw��8�Qc}�ÀI�(]ˬ����3Ǐ�v�
N���1	}.�O�����`����_��if]�"��S2p�+7�lݎ����1?��>D'����e8M �q����k8ҒGl�/s`a%De���O��0	��Ε�9�nv8IS:M�g�Njhv�v~�憚Z��d�c#��U��T���?�(�a��|-b�[����G�1w]�pR������P���ɐ����8�M�	Y�u��	� '׋�]II�Kmsx��j5DlJ�T0۴�YF�n���v}~����3�.q$N�C�[!��N��^�����T�[��M���sʏ��%�{���
��&��'+�}�l.���]��j��V�@�����V��<�F�1��XlxVHYEB    42ae    1110��!��BҠpK�	y�g��K�3������@ԝ[�q��E�Y��ɵ�bT9�Z(ۚ�=\ˈ�����f�\����~��+��X����N�6���S�z�zaG��`�˸�ˏ�� h���2�x��,�� �qQ���L]���i�	4�{r^�Q�5���V�O��_"���թt��{Ь_��X?R����d#Dx^u����򶌮�_��'V�İ�r	D�n��\��(�lqBxeZ:���سv����9����_u
��*e���0��E}H3	v�-
@?	Fk�,�D�JJ��촘�J�*c�Z��5�����'��Ӂ甽HL�A����i�f2��^�y�d/U�Y8����s
]�4
ӥV(6�U�[�F�06B��h�p�r�8�
��Cs|��+87*1��I m�Z#��X]i+K,kڠ?�N����C@���3��E@I��U�����D,0�p��x�3C)[4^�b�.��n�[�T8OF+	�`t���Ԡ7
�xZ�s4����C��{Ƃ�I�ǯ ���n,_�-�]y��Q��A�QEl�K�g�?�zc�g<j���-I:��]l��g}sGzu�<M�;��^�P�����bfPd�4d��X�W`�at^I�b~�J��BpW����=d�:>ly0TF}�¼�߫�R��BԈ�Y�#����z�S��C�%�!M+�����q�z�Z݈�����]��� 7�h��
�G�c%�ŰfE%�G=< �_�ݚ�����<�`A���⇒�m2�)�{΁V���UQ�7���P��'�w�����k�hr�ZmT�.��(T�P5��ళ���Ӣ�D�b!sB[b5)lU��g��J����S��)bN�����l���@�B�ƠDԿ���Vמ���{aa*3W6{�+�U�i#�t˟z�P�m95܋L�9���o�d,�|�c=�p�X
���7�;�3�#���j,�]��᝛�U��TvYhw �����Ұ�_�V�Yj���K�p0�����/�v�R�Rs�1_��F����Cڋ�^�
.`�/�u�[��4ȺpzĞw��3{�������;�~���T����7��7LѥD�I������<;�YJ7	v��L�鹻C�a3:�ํg�F*q��F�z��~t�V^/�S��
���0(�k�;^�+Af'4\�Z&	�ޅ��m�._�4����)4&F0<.����د��d4�T�p�;�����4����f(�r��ɕ�Cz\��{�H�VB���nY5,��ᒇ�ϊZ��.|�Cj�$�����"�sZn��g_s�)�iV��R�7�M�G�o�[j�̑u �C�*j`e=�ŭī.4�1���FV�$ۤ��4��Z�^C$Z(4��%o�]r��yR��R=S�￺n��L�|V�
���Ǩ�� 5�'�6���v|�(���!m2��j"���fu��|���D�i,�+F����ea�wy����������˙���DF�%�g�4��Xε�1��'\z�{�گ2Q�[���~ڷ\��-[U�'>!loem��R�ySq{Sa�b<�"$����Pp�яX�eV�'r �%{D�K�wA�߇n�y9̵�$]S3p�l��l�߽�)rp��{*����,}�e���_���x=s�>���p�����q���Z�E��j\��L�Ӣ��.�T��OH!\���������U�ړW�W������ϯ�K�aF��Ԥ�a��!�i������G2A��vk#��oE�̛ffGG%b�>M� wل�_A�)��D	b,;q�ǚ���ݻn�,�����YE~�+T� =zڵj]oe»Шyt��l�oNZ���ߓ�l}������h:�d@��y𱞆�P����b��⨜}�x�<6��O��/B���`\����<C�¦	��u �:͑���9���y��{�f�F�]�]����8L6�?&��^��X���
��t5���*�_Q	�il��N|��O1xSS��v�<D� ��-��X�b�0�w�w��匆=���uu����_S�x����ϺAn���9_���z[d��bCՠ,�&���/Ð�ط�#����A�ۣ�̎/��p�?�V:�K�0!�P$����#ߺ ��p��CG�-��'&��� K��<�����	=`�ˁ|w=�2���u��L˻��6�\��xK�\<=�1��M&���Ԯ��֧$~�؟1�޸���wI�C�K���1.p��~���V�:wd�D���A%��Ec=��h�q�?�-ie�0���S�d���,d����u�mQ�E[l$[�oMv�[�{��E�Rs�u���AƔPA��>O��:�?�D��z�i(�1*ǝ���Zn�����z��j3������MlvL0C���AA+x�Gч��l�$�r�/-�����k�>�f�*{�C�1k}I2�<��`SɇϚb���p&}=�鱄�����#s�K8���)��=n����� L��sp Ҹ��P�� 8���콿�=�����Am;��5���de\��^/~q?�ݳXUj�~W�iG�6>�!��Te�:S��S��:�����i�b]��<W��l��m���Дt���١l�T���Ȅ�)��0�`�~6Sg�u��AfqZ6UTHD��?�N��/�p�N�M^�0�WFED��=z-��`���$^�������|��5�������q,�����/>4�?:R��،�1����y[\�Ā�E9�&�T����|?�L�H�� j⳿��ۣO����#�!'�7�(?It��\�ݫ���%��m��� �� U�D�F�﮾��D?da�qc���»�J �q�C�䙫��+}�ĝ��L��6�q����4C�?������p�m\[]� �v���XۺC�g6ip���ܾ����� �$H�m�ruA�!��A�ĿW�x�Hm�<�
�����r�ws��ī�T3����P(袚���r&*�X�],�H�L�sP��dy���S*O&d:W��a�4~���Hv�[�jNy��b��A�9��u���s.k��M=��ę�ՕFs�)0��$OW���E!��q����-�#�r����nf����9�.��n0����MD���U�A��#r	'��&p�u�G�Z ���O�-������|�ZU���;�mBs�PzD���dNc�G9cGl΀S��W-F	Ƀը�.ϥ��<�	��J�s~���4F�}jL��I͒�9P��]���vÐ�A΍L|-��
�G�U-Wgf�����_���^^�6
�֮�n���ة"JaN�M�i�EU�e�a�p�S]f�&�������U��~��?�;3LWF�7�O��!5ZȼN�ed�t]��U��)Z�)$�I��-�Q�F©� ���o�ג�w��RS.�B��^]zL�� 	�T90�klM$=�(ss�<:^�a�-����k�B��3)N��$,ip���;�!6v.6H�M��Q
7zQ���fj �R��=Q5P�\��pQt{A\�j�	��A����?L�/[,���d�"���C�T���9zJ�$'��j��*�s��<�G���.��7, ֡������~EP�=m:x��a;���'����K�]�.��7C��F��Kc���;d*�4�`����X(v���#��\'?@8�u���i�{T���P,�-���mgm��=;�H�p�Bp� ��^���&�T*��{ DA-U�8O���_!��l}��'���8$��a�vQ䬮��.N|.�A��p�B|?�(Zp�myCS�=��[�߿���9>Щw�e�;f�E}���dJ�]�8�7�&v�ҭ=TZRuB�WO�ЏA���$�7�80�"����6��]��ڴ�I�v�����s�2�ߘ��b�٩�(�9}�>
Kp/R�0�	JU�����K�W���i�Vl=HJp���5���!E��?Ǚ�u��G������G���F�K��otz@vYi���^�=�?@	;bn(6� �K�f���0��˝T��.���6������`g��2oj)�fY`ń�\N^8��^��J�W����K1�J���*)�|�NJ$hO����]�>���oЧ,���s��T��ny\�Z�<聰�������},��J6���{��q~�+v9\iO�tTK�~Z8h���D�A�$� [�4M
m=a�h%�G��S#���Ep��\πCe�Z���&�I������+�A�