XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0�;Ej�MJ��h�Zqy���V�h9=�671����$�y�1�@M0�^�<����T
�3aϿ�ӽX��b����S0�k 5-��~�g��Ql�Nh(�E�`��`yZt�p(J�`��/4�<�}�ּ��.4����w�Z����^m"mTw�RrT��9U4��r��vnϬ�Գ�U�b��ct�\>4��ӣ+&ܡp��Thޮ�2��M  r���o+i�<�xM4l(2�.�z}r���Ȩ��:�]_P�7v,�v;]�li�(�C;x1���,��Ƀ׏ʒ������������>�,��5�0	�_�� ����Xr|�M��):&���D���jr���Ah�+Fӓz�R�N�[^6{,���]������t>��vFL�R��^��v�G60!���3����	fq^3-\M��9Q~k������봢�vL7�,��Es�x���I��d���G�A��p5@8��w����잒4�Dv�Ӧ����eI t�)f��|5f��I0�Ob�nW�T���������4��:��]�ufc��v�H ��|bg�>�����뽱��\��e룟ژ��l��[�D~�2?��T<����p9GoV�N�ob����#k����	�?�L_SE�9(�� �b����Qً�hP��̔�Ҝk����~#��@E�bì4���Y`�y�_��������^�d�1��Y)�.��P;S|�d�&RR�������������� �)q6��u�n���Ɠ�b��b?zk^]î &>�XlxVHYEB     f6d     6f0�TB��M�#"n8>w��r�]�8���G���pB��>A~�!ߛzd$��XX6�Z�]��ߝ�G�sU،� r�f�#�V�X�:�;.K"
�� � �0r��"U��>`x	ǧFB@�����J��ɲ�W-��TK*���\���43��U���e�z_�J+$:��x�^ki9YZ'a�n�E�6���z������>}oa��������x��P������Ѩ}Y���6�v/�8|���A�ͬ5��<��n�]$C�n��T@���Ǉf��_�i�,P=?Q q�$�-���Sp2�� ���'��1Љ��Xƌ{��ڄ�d��3oqt���p�d��p���+3�E����Y�%� 0�g�h�H�ǖ��蜏�6=?�hR~4�&5Y�PϮN�H�R�#��M�-T����^6Z��[�y�"�G1�8n�}��B��P�V"�� *p)4��q7X�(�m��ɫ�݂?�:��:l:ï�&�
��ןl)�	�^%դ��eؾ�!��qM��(3ǔ��F��v��N�8�[��)K#<�˵Ũ5�p�Sɑ��>�T��wE�@��4N�6l���EZa�l�9i��t6,�6Mmsf^���'w���&��/<ҪPY��ӠB�/����qT6��\��JO��X��ЪI��ʻ/�����~�l��0�X5�*~k�(����M��l�[)��C:ZN���A��=�Jά|r^c�FJ-�q�`���R����/�mm�41y������A�5�]��f�4��"��9���䓩�k���l�^g��T�
!R�����7��C����1\	@���\H�B���Neev�B�&�*[��UV) D��EM�7jdr�zKp*��虦��d���T���iN�ŔW��P�r_zxt�ތX�����k��, 
�҆}����G��VȓV��ʴe�voi�A����]�2!Yx�Wv����A�Y�K�"PVC�=�<�ծ���Ϝ	����!PCPc�转�w�\d�S�$A6:Lt���ȥhF;�[�ɼWT�xv#�U���,&��s�"p�{D�ͯ=�2Yy��@H�[�.hc��e�'�)�OlQDV
�۝�n����k��ǋ	+������#�`6m;�N33RiZ�4j<�P���s���l-heS8�i6���Ӝ��b�����$p�D���ٻl�.g��LHN�����T^�:��¢<��(�$=F�޹ab�`��:�t�lYO��~��E1+���]}o�1��-��(Lg³(*�r�7����Zzy۾�H;�q�I��I���S���G��M����f�y�]�kf�G���&[�l��k��=r3d�t��k*w4n�XW>��
,"xDc���m�#u�ż:Y��{7�y��{���Fd#���x�AhQ"�|YuR�Ȋk����eD�w�]�c4Qt�٪۠k�YJ%�	����ł��[eO��˝ՎcC�e>_}蚶emFS? ���O�Q�w���2iw�q��bA�X~���N�:q4��"�^��^��{�̰�b�	��q����w�rk�G3�ɴ�8��)�\��[阯F��J��#���ڵa�|I��w'���!\�L��l�dߕ�SX�Ϫ�c��&p�3i\��2krl�=�����jh��?�b[ԍ�!/΍�������8�2���^@Y�GB~=5'F�XPnv˧s&�����s��ն���`3��[��*�
*0|1�� �YAs'�Yr'�m�����