XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��=��zn+���Do�܊g>D��&%:���dS�I�Խ�����;�X_���PS�SSU�(��w*���79��b�('1V����N�(���H*����,�y�K��wm�����{�����	s�Ș'LT����T���BX]Kx1��Wts�k02F�E�)Ly����mu��`(�$�?l����=h��UXх����t��H����sD=f��ĝ�!�9;IE�����]����L�C[ �Jպ�S��-�����Z
�{xn��)Hfm6-��J��!���F	0	�͐�ة;�gt��mk�Ol��&�'�YI����Q(��"03���oI!�lM�}�%*NL�p�˅G�
w:�9�1�1������ND(��n�W~Y!�Ia��)f����u�����/�[yǟ�|���a��͢�X��9	Yd?�OY�yz_kEX8�~�a|�^��u��?>�[���4fM09�Y��5�8��: ��Lm�v����.���V!2Vq$��0�/�-.H�SL����+�+ uI��.L`*�l�,'���^�'ogbL[�ki-��0�S�u3��.��G_l��A+����ےE�����S�Q��S�8�>�"0!F���Iy�%E`�l �Id
g1�(Y$�]%�MV�b�f^�8�w
08� ���`y����^��Ƚ�JOF��(�sc�,�-�`���T�R�O�P�q���Cg���܆������aV8�9��~�Ҧ���XlxVHYEB    3b09     f80�K�������df��*0�ߨ�R����ɠ\�OnRY��Ob���1/�5C��^��w�ǃG2*�!n��u�Gz4$&��#�f�qf#���y��o��3��Й�q�����M�BQX�P(�#I=Q���ęL.=NE��]���[��=Ne��2\o3�IH#���E!_��{����E��Ǜɵ����W350&���@���^k͌��콑W4C�7[d�͠t?V��?���N��3�Q�Un|oI�n*�'dx+���d�ӵ�h7�D-:���8�_ W��=@D8|^3e�?k���!���jk1�S.�0��M�4���I')�'	�{�S�v�in�4W�ʜ��U��=�j`�e9�0�Ѩ%��ݴ�Z�g9��ڙ�P/�(�r����D���aE��݉1��M	א��^	�B#��Et�&s10R��18-�|���S&/�]��Ts�+�������)�lP��2d釘�Ngή�����eD+���T3�b�f��f/�H�
�w�0bz�q�/چ�����g4ǭ}y�G�����|J۶|���:�����t�U2�F�b��s���E�|t�y'���H�p_�8]����3����q}*$�]��c���V}�{�e�jw�f",�+xT�@_	lah�(���`����w�Z���	!���x1?+�>Vuf,K�Q(̙T��V9$�����t�T�(��	⇁��H�6��'t%�8s���hW 97��("f�0�)3/���C����"Px0�0o�=���ٮ܍��8z٬c�բ��vޟ2�G�c$
�3�-J�����3��!��l�o��^@�62z��E���2~���%����O2�h�,�3*�bFN'z}�B�����f-ki@�0�
�o���9찲q�!jt��S�)�L6u��_����ũ*�z��HqI��oK���a'({��rK5�������a	0Gf¬-�a������g^`�|N˃n��e��g��M�B]�/��a^,��\/�`�C]sB#[s��G"	��y@3�V���隶��Z�$N�P���>��d�|�&���*t�7���cifO�?'m�����?N��x/h˂l
A�*��	��3�m�f���V��0)�M�A��Dw��u�g�;�yW��\��x����3Ҙ5���xc5�ܿف�	'�o���lW\J����A^���p����V�1�ʹ�=��<�\7��KY*���f<C���H����É��*���B?���Y�s����<���)�O� a�=����r�$�*vnT��]����=���?�d�V�X�����{�G��,K,@1��O�!<�6�2��0�wUjC^����D���iOku��(�?,�u�j<	r�a9lo�g��A;M��Q��y�[���Tन�����a���.�8��|o=�C�te|���y�W.&W��4��hY��V���i��#j�k,52%�kJ �K��0�uft(X� ����\F	��T��1c�Qr����5��@�F^�;����)n�x	찅����̨����� -��6�7��P���H���k�"2�YJˇ2��E'R�h�7��s:�ʳ辞_�����*`g6�zW���B�~G�4�����r�e-6j
�RP_�z��e����1l�w�k:�+7�2�-����ĩνܔ��q�|!0W~Z6��r�l���
eÃ�Ge�0��n��/�%�rt�:��0v�(a�����.
���\p�- ��A�PzP�\�n}�X,��*���h�{�l�׼?w0[����0^�����%���ڒ�����\Mg���.a��6���� ���+S"8dc�g���G��0�/U{R�q�g��g;Z��4L����yo��������pw��BیՎ��t��"Ɓ`=`E��f���y�V
�/��M��,[۸��x�W������G(�m�y�J5�!(��������s">�zH��{�8ܢ�G������P��6r׸j�P����"Xa��x9�n�g!��H�Ƶ{	�-yZ�}�_v������5zbC�$��jn�<�y�p}֕��ߗU���z��8N��rEq��"17.���Tu���|�N�5`Ǳ�ʗ��m-�/�����C�A�ei����W�ڑ�ة���.���Q`��z�]K��mi�'�`X
2Z�ő�u��=�<�\�b�[���Dt�m�rV!+����#��%���H��;WT|�z K�T�eD�/�ҫ���gŗ�<�����J���(,�_��9���$-
�3������8 �*x�
�'��}���~LEK��n����}�'h?�~��\�1�a^6٠���w�?���N渟��Ѓ#�k��x�~��,�%��qQ�J�YŹ<�MM��l2����u�2�Č��8f҆���oy�P~	S�����'3���À$L̶L{��'��s�N��f�� ���GM�k`W�5��F˄|��z����%̅��x�����%��j��b5�-��r�c�<Ksd��3Q������:������j}���P	�ݒ�&?Њ\�Z:�������Zӕս���"�V;��8Z�[�h�Ŝ%H�③��U9���A�&Ω]�He�)j����Q-�m�N��T���߬�2:N��É���<��t>��``w"A��$zm3ϳ�^!�y
ʃ}�5�
�����;[5�b�$,=�~�K�s#�Ѣ�s>Ϥ�����d&{_NZ�{�y����J�G|v9�p�ΊZΤ��ִ�Y�P�V.]�d��weQ�ە�t����7�ҷ�
Ͳ[Ո- HJ�v����$~�gZ�"�pϦ����/�q�Q�,T6z���Yn�q���課[��֨&�?(&��v̠K=w�ˤ3+\ȳ��x>�J6��R���D߉ݴϠ�>�%_ SL��W���ͣI	1�]���,O�ck �����/����gz5C���g���,?�Z=?�W��,S��k���:�ٮ�i}}��i�lp[��b'��w2�Am�rk��۲�� ��VwIJ�9���t�
�8}�R�ȹ�i�|3"�P����9%\�^;:�څ���2V�����M����#|�FH�	�>ic���7�ąW�q3�ܓ���/4���: H�j�X�M�C�����=[��Wë�u�C*i^n9�#o������]7�=����LE�M��S�����X��^�h
��~�I�G��]�b�9��zÁݝ)�\���S���u�����zUsW���H�7@_�����d���q!^]�r������&K��Z]�a���r1X�U
���|��?���h������U0�O2,EB��N���W�&���C�p��@��e�]�j`(@�D*4	k��M�~�q0�Tc��MAF�S�Q=����5 �Sf�AL H?��p������&�XoF KФ�}��$s߶��)
Z ɀ��+L;�J��Zk�]�#�%�&�$r���Ck�+��]ꛀ���N�Y_�tYL�7�����$�ҟ�ߟa.�	'i���©6�I�/��	g��Z�^�Q'��?D�Ԓ����9f-~6����X�T�!����=�Wȏ��a2M���.���<�R�[7<wwD�����9�|G��(�S̓:/M4/�Y��"On�+=+X�_l{�X g����?!c��v�`�3q�Y=~�ys�,��!5����C#]���5�O%Li,YB��H9�(�iа"nn�M���o4�7�jм/&�#P7ҟ���3t����:����rUËs�*����lȶ�[�!��B��b�ox=�],k��qV�ԃ�)o�y�u0r#