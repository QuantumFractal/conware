XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���'�+a/��КBs�U�8�y�����S)�}wF�;�K)�}�m���!��$�,��G���l��=��ITY��|�N�eBY�yj�����9d��\l|�U{e�1ůB9R�̎��l��[nɮ�?�L���c�6�qJ���ŗ�'�+�<�Ve��N���I]��l�����e�Y?	� sezAz�ǰ��=n(c�C>T�1�-��<���k0`��c.�'�	:�HZj$�T꯬�oli�V~�U��-}D]K6z#E��X�f�<���X�����^z9d��z.��+��kОW�1�w�H ��U�V|�]P0�e`�ɞYΥ:0i�<&�D	��օ�4jR����n�����xT��Yj�7V� 7J��[�}p���6Ƭ��^ۀ�h�jg0f�AY��k'z��N;L*�t�!�����cK4�E\F7�R��*E4��d&X���~w��䌓y��QM��c��Gd�����0���(v2�r_w�Y=:��u�6��;���B,"[�d�9�$�'T����i�vN�����$b0�Y~|�A���7B	����\B0�bj��kT�:�̹��^<���mz�N��v_���I�u�~�%�����Q��3F2 ��V]�O��(,�+�̘��Rә|��l�x;?����ޕ��fW/��]�zb%ɂM�__����	Ǻ+���߁1Ol���V@����M��W�v�r�k�Hծ�̩@8@ Y�҈Xvw����%��D�(7�"��tc�~��nsXlxVHYEB    42ae    1110MDGSCn�h;�?=ܧ%�� U�7B���-bb��b9\�B4����������J���'Wʋ�=pY�����4� DL��+�R%ϸ�l�d�� �c�y_[���g��d��\�t�yd�>[=0��yj�|�=xw���v�iگ�(J�vm�]6�1�J_�IHZ���� 5��=ª~ʺ�H>3�;��kL~��D)u�b�ם"����F�:�� �6}�	��hvb�,�$p�����/�c4)��-ɿ�ES����̟$鲗g�ɼZ�8��6����b��:��Gbz&�3ѫ�H�!d�2Z#:׳����aj�s�w+�i���G���K�m�K���7���A�@WpEE����c��
�!٫ 3 �PE�՜��y'����O�U�	��Ђ�d$�������V#�P�)�7�O��4��-��m���� d�pN<�9�q�x��#�X��
`�M��r�a��M��2~B����8�j*l�iLՁ�2p�6LcF1�6x�+Nh�+�*�֞
��bA��Xg��fV9o��y��M0�8�m�u�ۇW�lr��qCʏ8���ٱ�-&�4��R�ch=U�7�Y��S��NɚD[W˱��݄*05�����)mya�v����QG��ts+߉�XuT�ʁi+ǆcj���!l_��
-"�ɗ�Ǧ�3�m	�]�i��}��'��+}B-C59�L��!�`很���9�j�B�O�T��+&RH15	�DG�
4TD���P�#>	����B��"����_�]�r��a� �IQW��o\��S�-�?��L�\a�ʻa�b�����Z#��킆=/b�(����-i/<����Df����g��w��\��:/ �W�ns�f�ҡn��p����
��vQ�]>�sO�����);Vؠl�e@��AY�8��UU���Q	KT�k [��8�.����Yz���.��^)ڟ�Q��sx�����7�`J�2��˛�C���;Zq?�R��eLptυɁ��*�_Kd�Qn4�+���� 	�HS��P��ܵ��#N0u�q_%P
��/��¢��7X���n,@)GtS�C;��,w����
Y���{�Ԃ�|ֶ��/\�L<`j�2�L ���₱��̯צl�x�#Ct;R|[��T&���d���Kmε�H����]��%�m�ظ�b���
⽉@DA���`�\�p�W@��PϜ�	k^XI`���U�~Z��ce��MԤi@��{AMQ5B���sVMH�YBcy;�����>�t��빦�]Pf�\�4Յ.8~/�5��ւ���E"��G
G���@��rؑ�{�F�j���Eђ�E�t���*ņ��IJ��O��Y]O�_��uQ��xC�b1������j��/�$wi���PnG{�ް�>��Gb���8g�=z�tμ���6�|���X�ꀽ�W���_� ������Ŧ
���i7��X_��hh)�4��'�3�����F�р�lӄT��.��+ɪ��� W�na����o��b�r�4�g�4����n�)�؈��:�Ɏ�/��?`]����^Hx�0���/j��"�Xo�x���{���75q��EIa��8�EQ�+
�-��9}{Y��ֈDP��65ҫ��߾�%FF�_ǹ:r#��MjX��W��Av$^	m���Nɽ�����8��G�֠�8L�1�-�;$"ؘ4������:���q��<�����Z)�&�8q��r,���L�!�F�xc�ΕܲM�E�!!�f�_��a���E�|/*m��Xu: �;��Eϖ�'>�a#�k��@#�DT����Y��~���9@�\��^OO
jl��n��|G�0��{h��s�'�<�I���wɠ }A�;����d����ܱ>&ݭ����M�&��Q��ʐ0�+K��x:Z�\c�[�֑����V�����'8^�����%�b�L�Zc�I|+�r�j�:����a��h^V����̅5]u�횡^?<����g�η(^�PP^[Um�#�CＥ9h���E�Z���rn")k�u��N�����J��Dt][���TKqy�O�b��ܱ�G������wc���3�=$�A��dgWD�E��`$��x.E�#�=yW>/,�X�L��Q�(�V)�ĒR<�L5k�׬�n����H,X�I��]�=>�-�(-f^���)�ʅ�C=�І�|Yg���ՙ Fl�!�l�v�)ŧ!�;��o:Z����H;�e�3���%��e�T8 ���#n��>)z����"�cVt�w8�qJ�:��P��@�敫X.�,�i8���+	��>����꬇�(�O{�U�������KW�%�D�����v��� 1zr�mHʻ�����;:Q^%4�>��w���1t��m����*�ť}2�(ߣA�),��#�(1Q{��b���w+%+���P�հ�U�9��X�!s3�2|t��o�F���D� ����K^�5�zb9��%&�N
�4�[�YCS�|)X@kB�J�,5�0U���8�F�.�p���=)�R�w �%�u%��f'φ�!������K�(v���|�����MG��q[�?ن��|�_�m�x�C����+Eg�G� �6YNk`�7Fה�FG���p�������g�8L˦I�O0�q�`N.$6� ��&��S��kؘ�Gcg9���1쁛K� I��� =��w25��m���m�ܙ�D���x٩s5b�p�B�r�~�o���!�ۃ�F	¯n���O�w��]�h�|�۳ڗ��2`��M�r	�j#�*���~42�Dz�����z�$S��uqT�t�p�_�ю��W��{����u�G�}���m�lb< ����|ɬ"�ۋ���]��8��!�K�v��"�6�����c�{�0����P�$	�`�⏻v̧bx�@:¦����G_q:v;� ��\U�8	7�݋��t��gci�r28L��x Bi�����f�ڔ��O2�#Qm.�Q(�=���ԙ!띜E�M3��Z`���$o����?����*Q��}�?Q-��l%�=�qK�=��2���؋�O1���9��脈����3���w��#k�G�,r]j���������!��ۃ10�8X\٨���=���H׌�+6�@U���1 h��B�0��{�$��H����n#��'v
�FB�J&������p�� �1h�`�����ܦ+Iܼ�.�;�7ka9k������"��}�]�X�@�_3������!}k#��u1�>]�V�=R��!����]��R�b-pR,�)�H�X�)s���a	�)� .�,�L~Va��SI�x�운@'�������3�SIb�P����������Y	?��(�Bh���4첁�k��tWVV^2)V�o����D0�E�jdn{h����6I�.QC+��E�}�xKJL�y���M�{i�`�]������>�ʽ,+�"Ԙ'�!��
��v~�m-c��#��j$Q�=�#.
j����R�9��sH��o�y�`�k�[�}_bN��iw��!�1yA|�[t�
U��q%�v����L��uІcB!W���Z`�~�yX� b1R�+��kX�:
*7o*��p����O=�U��Г����8`�y�+T��XHQ��1�(�{�'ԋ��ﺔ�+b% *	��ݤ�N�v�E�[GuJz��i�:%(�� `�Q0�ŀ�@�O�ۛ^ׯU�х�b;T.8z$b*C������u�"��|�@5+k��ީ	�&� ��}~+Ah�� ���R�Z�ŎA&�Z⺑�l�G~��l��w�ޞ�o)x�Ƙ��k�p���Sd�!)��cSK+�IT/�?�c��8$~E���BS�{�:���V�*�����]�a;� B5 �����M"�j$�.�����@��Z����7���+��	PL`T!�/]�M,���QY�擻uuS����?R��
���K==e� Q��U���s���Koű�<���J�y�G���ӣƘ��E�k']A���&Nc�=�G��Q���(�v����&-#�eg��@�t�*���L)J)�N�n,'�J�\W��w����Vd�5
}����B4vW�w�Ǽ��wf�`��WW	ĤY/����������I�����y�1�͡�9��:e�K�3h{�+��(��y԰W�/�T����{@pn���14U�E�WT��E�� �����Ӕ��4e�P޽�l���ܿ��\x�����N�g�j$�
�z���q29�W�_����5��F�$S�?��(N����`m;<�.�J���I^ 'u�e