XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Y�9��<g�x6@�ܩQw�!C�
y�I~�XU�T6[��Z���`��۟8�Qt�";Czpz�ER�=�E���B�a��^�sXR��[�\,�THrH��H1�)�;�>dr�Y��ԃ� �k���@0�M����;(���nq�"1�,����Ꭼ]��[k^ǵ���!=43_��-d�	���a(de Z��=�)(6��A�F|M�o�����'��5QՒ3 �v��^��uOQ���[�ZGR�8��f��e���*	�:���7��r�z���Z���Ƭ�M��G�z�C�F��?i�`�AN�U
ߠq��4]03���ŋ�ӌ,^�H�|�����Ј��`�����u�r�����%�0'�F��F���������p�*Ssh7˖4� �J�1����Q�q�S�</�Ĥ}3��)U�5ϕ^�R��lށ
��7C}�ߗo��y�TG��Kx�1)��_u�uƤ���l�{F�����!�V9�ѽ�N\��8l��|�����w/�Fh�`���!D�\g�pP�
	�)�k�# Ti��|M�ݰƓ�AA��i�8NQ*rZ`�|��>$��8�{wx
��'u��tR��� ��+���X���>x�vE��=�����z�gVku�>d�x���{O�Ə�#�|�@�,ge�Yߴ��iΌ
�!G`��Vo��oƩ����6�[�5�h⍿�0ps�y:��Y��.�`C�.��{J�UC�W�C�]WP8B���ݍ������dF�H5��]M�XlxVHYEB    b3c6    25b0W��`u�p���;Vs� p�?j���!��q���ֳ�\�֥f��&��ḳnݶ��鐔��:WJ�M��Õ�.2(��Y�:�&�{7yQ'�=�ӸO��1��٣����akZT�\Ω&����󈥃Kl���4�wwa������=: �X�
1���!��M���)�/@q�S��S���3"��o�5�S�~�ZƩy��#�fYV0(�88Uɑm��1�Nu@����|B�{>���פ������?�F~!�v/�N��dr�?Ԋ1!~SjrH(�$�E�D;5�d�85}���u�t\����j=� 
�F@��f�	Ҽ���Ĺy$o;�Y�e���,)q㑩'z��=ܮm����:qr�O"#���Ɩ�.��n#�
���4$?�埢�U��Vc�V
��c�$}ΐ�;U���讠�s�f�9�r�|�r��h���򃂫�pM���H{6;.��=yW*͟k �7c%_�<2�M����!���}�笉��s+m鲩�4&�|Q`O��w�":>I{Rj��t�]��Ţ�+[dۙ�z�2��$,�ѱ9^ཋt�l��#��! �,�7^`�W�IZ��2cC*B������3��.���L��P�~�I)�px��>:Ձ��ځ�$���d8<M�`)3䠙�<���L�c��W�_D�V�5g 6�V��nP�xf������>HB��Ϟ� ,�v������uU�J�&aZ��*�R�^�A	˳L9/�؎���Y���ʃ��Hu	`\�+�g��K�Y%��WvBZ�Bp.[�Bl����b���%�?|$E;�}b�Q�q�xQ��J��<>%c�z�0� ���ֽA3�
�nA�P� "�7Z	eH�
���~��]�����oZ��Z�A!:���˖�[�&�!Q��MG�W��� �s�P�,��� ��9G�.q �`N��?^Ă�2{�{bu�?V�@�����j-E�	��6f;k��X��7��7I�[FE���/oe�>�/��侬P�;aZ�.,ug�<�E�⅌n�©/$S,T��x���Y��|݉���_
�>3�\pԕ�B)ϧ򪾬��K�y�+olT��t�^���,�W�}�gL�c��K:��l>�#0�%�N_���q[���	�6әV��Y� ��J�2�6{3�2p?��e`w�5:Eߍ�w��7��O����.��J�R��'����B�Ѧ�${�#�|�T%�̅H�G��&�L�������zaa~����Єh�U	A!���`��3C�V�8l-T� � I�ki�ai(�L�'#w�A�!Ų��	S*��}mі�b\Rbg��u��:��S�(7��z)4n����%kuɽp�V
����Kȟ%��s��2T;�AL�r�½CK�b3�L8Re���ӮN�l=+3У�����s��#�����zsĤ��XԒ���]r���'�mL6������!����~�V�}K�-j\H����_�Z|�Ҹ���R%�0�y��<��J���kA/S/��� �)|�Zat�t'��s�hB��B_)�G?���,�V� 8~��1���CE�?L7�W�$RI��mfj1H�]f����D*X��<�3TH�f���|������3�5�g}sAhai���\0[�th��q9:?��j:'��̜�LA���+�|�&���3b�B��#��ⲭ��#�7g�d�҈���� ��(އz6r��
�|j`��(��E�X��N�顬o�="�?�����8�����m��i���Cj��Z����h�~ RWR��2s���I�J'�GN6���f�B��T,�޳�	�W;��j9���"t����%��(zN,%�O��������ӣ�JC��P�1��C4MӤ���V2K��a���)l>��|�)�6�/V0h�R&�� H�Yh��W�q�a܏r��!����.�ZW,�e.��/#�p�Ǎ���Ůca�2�ԍB�a�yx>�M�*�E�=�r������F��,��|=��H�F8��+������j��Ġ.��+�t�V1o�O8ni�C���|+�.��Q��T�#A$�}4*K�v����{)30��=�1.d��cPm8!1�M����YY$�����Xt��B���`�|H��%:T��2ˈP@8���y?quJ*�	X�2����*6ZTՀV� p܏#���
N�tf����P�.���\���g���/�ҦO:��:�C��AIR.�/��u`G���K�k��Wm�Z<e����N���?x�9TO��6�� O�%7iT�/Y�w�]ʩ,��я����B�;�8U�r{��Sfb�)�y;�@����
��D�mUt�MKm�g�$U=Y���P��|�Z��=�?��v�L#w#���:A��'��Ѐ��%�OB�%�&Dr�t��~�������- �r�u]f�s�]�C[���:�Y�c32C����F�t9��A��(_��m�Jv;�+~�s�Hʑ��y=^	In���(�ĥ�_��m�gQ4i:M�yaX���"ά���Qf2����-���$�I*d�\�����a�f����/���9.�dZC�bei}�<	"b}-X�d`d0ߒ@\���ѝlO���=�-,Q{���NJD����Nv�q��[gC��0(:��_�������}�.i�p���浘��c�1��CMGD�*¢GD�dϥy��nq��_i؟*�_�jh�1�ڋ��#>�9
�ڦP9R�^Mh�p\�̭H&���r>��xA}"�"����� ׶)�E�0�0چ��'�VO�	�+a������-dǤ�C�v�8?q}�()��F1�����2�x���-�7v��Φu��yg�j��!�P�l]&-�Dg��p>����T�	Z�D��'I�S�����zM��f�����G�s�r��3����f&B��t:���qW\�H�-g������y�>ᇡ-� ���;�����ω��y3ְ�e�w��r����u�uk�(�v�'U�G~g=����>�Q�$���$=��i�IF��zx�����j��{g�h�*x�:�}K�0�f��|�*��rQ�mm�ƪ7-�����8�Q9��m-��r�<��]����_xT���['WOˤ��0e�⭾��ٟ9�m��=LyxO(W͠*��� =|g��m�����&m%�-G$ a���zu��V�S�	�吚ht���Z�'��4*k���f/!7E�ְ�k*v@r�X��Y�N�hQ�Đ�k_�\�������0 J���9�^'��,5;�K��z��rwR���%c�.O�����9r���V�CòM���l��I��V{����_F�š*:�r����>�(#9�@;�e{C��oIŶ.oȽ[]��Ƙ��}i;�$�q�rh=RW�?!t��K�p�1�;��|��XJv-hTV�n]=��a�r��{����_�{B��2S3�28۞0R���Nv�+������w����P�?.|���t4_��]!��;�֫~>sS���G$]~��ɚ�#jZ��,/�����:'�mx���*�k'i��v~땎+?��oTGQ�t��&�� �լÌ�	|�\�c�>NC�*�岓�a�+0B|��7)@� N�'2O�����������zA9�Y���dϝsW�!�'����=�Wk�IeB�+r�5/E9�{  �a)J�x����vA��� O�W��v������ɧ��!�`�k�	���3u�0� �-z\�����#�s���S�4<���;��W��}�8�|{�pȝ��_y.���[�~�Ma�Ci����v{D#���ë�����J2������^�����6j��`�9��
[BގX�FLFQ�3`�<�fKs�*�\�ĵ��L0�_a ��i���-D�F�(����~���V\�� �HƿBg&������|~�TJ yQ�
Z�#�&�Fȯ�S屇5�d�+��;䀫��P�[7��J]~Q7LTA���>����=� �=xv[1���3�j��1���8�a�
�e�>+g��v�=X��G�x�ގ��&�sl[��|�j�LN�1,/�{���R�N����g���f��)�;U:���?�Uĝh��˿g�������7<��'��Q�51-5�5IzJ�	b�&=�t-⸧u���M^�L���@	v��ڙ�E��e�?�K��qz�����kB8���K ,�EmI��I�:vӜ�l��C����}��[��̑�,�*K\�M�ܥ���ߐz�d0fſU��>N��@H��Z����9l�y m�9nob�=��|ez�EޖL����	1�8�ε^��L��ʮ`ޑ$��4Ԁ����M����MQ�ݨB��;�*�,�"o�>�#$)0}k�eB+�f|��1�!�:6�яڣ����ǘ�"� @��b<Hm\����$r�į��V�F�j��=�Tko�<���2�pX��l1*C{���@��٫���w"��2�YS�I.��*��sm��-(Oq����~-Η�SΊ$p��7'����I��TA"'�X��N�-Äu���,�)�VL����8fX�YTW.���拔\8���r�tZ�ȸ#\ �%,)������%�S��� C[�y�\9��豚W�o԰�������j�����#�E��v}��
2�G��nY>��Q�(����o��|`Ao���KCN�=Rv�ޕ�����o��,�)��:5lr�
 ��.#'/��՝�;f�P���Ħ�lT,R<�a�J!Fq�E-\�i{��ۣ٤��I;�,Q�,�ͷb�6Ǹ�a�ס�i��8��(6��qP{�^"�CW��+�Ф�ȪP)A?��W/A�'��x�Ԋ��6�p3/��������<|�����Ż���<"�_,����*���?�mo��>B��7���"����D����%)��E���L�{�AMͣ�� ��̌k������uK�h�_�ks8���C y���a*֬vՓ����fξ�i9��q`�@�j����y����_��
��8�$�`	(l�r5�zfZ%h�	'�� ���"�Y��>�Q��u�/Co��$N0.� ����[��~[XU�Y�*���|��L�>�r��W$�IBOF#u ��*hs�)�!'X������I��ⳝ�$KG��G�k���&�~.�Ax�������f�����rɢ}}
� ��F͡JzCf��}t�g_+\a���b�q�+�cꀹr�?b��;�oc7��0��N�M��@M�Ѩ���G��Y����_
�z5��}��
Q�L�vF�j(��
p���+��L�|�8tHD5�*��r�M����t�x�G�P+��\E��e���e�М��#�����w�A�ݞKiY�����\,HA���P,��J-q�~+��nS�auqîBK�o�<N�	狶�B�f	��v!"\�;��O�9�~lFI��=�lr�M[��jc� I�n�٣-�*&!��L���82 ��>;�Wv#�z�u�^��r�gO�����������m����c�'h�o!epQ���*剁s�ؐ�8I�,����]� R��7}�z�{�*ǰɾ$͐�,62q-���7N�#�4%aZ,/��>�6�ձ�@����Vc�!����lŎ(��O��g��o5}^�w�n!+���t/%�|��Eե�Y���hk7t��<��TK=Q>����9�
M_8
bb\=��}r\��v����7{n��[Y�w$4Jλq��E�6�o����ÿ�qQO����+J#��#|;~K��O�ݦR�7�{����*�e�~���Y��1�?mY�w�i��yR	<����*��K�zZI �0�t�m��h��K��]�s�V�D�=�h�������嫽>g����T:=�V|��?�{R��V�����u���*l���~�P��g�?߲GVd�*�	��v<�K>u,~�H�����M��x-6��� ���o��֚� o��+��2�VK�0��ۈ�2�F���q� �9�b~�m��I�j�g��P�Fj�,���P�ǹmoܘ�sK;�'VSҍ�f�8�*C��܏I�\�t�Y7�+� �;�$�r��k�.��Z���(F�ۗ],��L؂��;K���*<%�@M���p��8V֩{EՌB ^o\�8s��f���ϱ�MY�KC��9����{|�l1��y@���8s��1���]o/g�a��^{��!n�����fnj��yW���J�|
��C��Ax60/K@�����t(���f��&/+#��H��� �� �f�!/㝸��|��Q�۴z�8�]cPH���Df�z*w��*.g��i	�!i�2l�g��-^���i�tS�7mckƱ�3$�[��0cEKw��B�sƔ���S�b��,��H�92:�/_����)��_�������*��R6X ��dT�7�;��Z/��kå�"��-�X(���Z�^2��R�[��L�ѱ��6t�Q*\v�]\y���`}\7�͙k�W��� ��������;�������s�!o���u���-o�z&�r�������G=[�n�Z�=�ҥ����Z�����#/g��?|\a��� `����Q�W�A�>��_oQ�=�W�oD��sK���M"����C1�(������<�2:y�?�����o�FS��0�iz�l�6�R�v4�{/����� y'g�=)��"±mz�Rh�$�#uv����N����Mwģ�%��r�Bp9� K�K�O���A��,IV��.�F~n�BP܁���_�'O��aCyB��rw��e��.w<}����bl�#Dil|��o�F��ŝ�Q�\�U�͙<Oq�v ����L���ͩ�����=���~ ����voZ�>�Z-�jԩĎ�[�WA[S�&dТ�G�n�R�V7ěe���PH�C�K������`��(�Eϔ��-��R�L]����a�x>����^��!������EG��p~�1����0<͉��b"M}�Ol�Z̓���ڞH�f�����9�\�	s�9k!���Q�v|��J&�^�������{v�l��Co���G�»wC�������Wxgh�G����*T����f�q{�`)D
7���vπ-�S4CFx�Z+;�șY L>��#� ��ǔ��&]ONv�Q���ً,7UвQ�
���A(5�Y�x*�b|k�Ȟ���������yͽ�J���Me5!��f���}�M��g]@�ƴ��g��͌�Z�i���۲�༪m � Tά)����	���<��խ���(�����L����Y<C��γ��	���}!tm@9�����^]�h B.m��l�ö1���]42��cI&������a���/��eӌRV����F��jú�D.�U������(g�j|v"�/N��-2��0����]�����pJ�5�W���|�lJ���#�L�ae�����TB�1D�e���
S*��o>�`Bi��ΔD�;��N����ܐ]�{�����t��/WY��7��fR�ɱ	Ky��[����+y��>5	�Cj)8I�j8��%\Nc�'T<,��]�8��ءRi�km�*ZK_5Q:���5�C�F�8�v�`��x��O~�-#�.���Hgi���Z��S�Yv�Cu|������<<V@�,7]�3g`>b  �f���Aj�\�曉7�X�^����B�!�(���bn+�Vk�-[}X�[yF(�^��le���	Mn8<!�M}�~�R6�2��ت`���*&�b�0J�g�"Y3���x����p�̐�ȳSf��*�X�~������4��H�U]���#�qsT���*��@T>�m�+���e���t�B����$ï�}wE����;%>��e�ΰ�B��o��/�o�5I�G�b�_�a�P�qI�?�E+W�q�R(���r���j1�tߪ��G��/	�[5c��Cp�k(�ą�N� k@��s	�jtr)�Vy՟�(6��w.�߻��^QJ�(���f�iz��A|�r��#������6Ë)>x����ӴjgV~/�/vb"�^y�\���'� �ޓ��4MT��r�6.��l�mn}����g0�MéD1����z��u�T�mq�]2�ߤ��I[�M�U��΀���q��U��c(��=�u�-��A �v=bH�Z�����tb���2��T�p��I�XD~��*�w�iؘ�.h��f� dt�u�/��~�ܥ��ی�Xls��Ó��j���.�aNF&w�������B�(�@��i���8��(������sV����"�P`d�|;/���@*�ٓ!iN��p3��r���}��
n�hkCL�Ћ�VN�f\d�"�mi�N��ϣ�IY�6T��!����'o��t�����"������������s�K���:�8�E�����p-8ۑ�`��:�>�s���'�i�9Z�^�\��@���(!`v��1��#^�Q5;�L(�3xѰ�:p2V�M� ��V�/e���O)�RR�F�����H�|�$����+ѹp���z4�d��8��p�����w2K��&��\zK)����W���u��[���Z��
��z+v�f���wX Ǒ	{`΋��Y�]6%'I�2�D}G��u���y��l�B��Fu�N&?ԖN@�M��2h��Whz���#2��+H���pW�w���}�P�b�3���	[�B4Č�G���0dU
�.,2!Qv)�x� ����8-k��y[�JSP�}�a�V����=�K�K��BR<��mEJ[�r�W�m������sb�	�<#����v�T
ߊ�^(r��)}���|Kt�D�(���@���K�g|Խ�� �\�y�/��@�x>}��"�t�19T\KU��bYe=�R�"�sO2XS6/�`�( $�q,�"߸zguH�f������0ܜ���7v���f���8��}�sM��E���sE�⍟h1��y���l�������H���J14�Y�i�L�	bn��~��GTs�p�߬�y�l���M> �4��l�����u����vֲF�˶�=>т����&Iu����er/-�?	��7��]`Z~A�~���j;Q��4�_�WXg�3W`^VB��w��j��a��5k��͎��^�G��7��@��BD��ä�rKrK�Y��k�� �@@e���ƃX���PlsG5@o�����O�&=hǱ@M�g8�[�}�h�$H����6�)准F���8i�J��'�����؟<Z�I	=���zn�i���x����b���S*>p!<SF�j�vv̝�xoє������Q��V˘���l�9���x�S��� ��P-���T\�
����8ʪƴ��<�x?�ճJ��CE�� �y�x�*+�y�G�_������ RGk��6\m�T��W�[1Pb}�RB���?�sh�ш�p