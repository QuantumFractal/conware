XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��l?�����l��$�l�.E8[(P���֭X��;�NC�c2@~X�(��\���?��ƞ���=Ȃ��,�(X �b� ��Pf�W(�v�X����&\��Ě/��4I �mz7��S�G)&���=���zV�
��o� �Z-4�{#�7�֎������hF�k�tռ��&�.��S+��e$L=#�oa�S�rQ��4#+�pv]���]�HR�`�N����|w���9�R�����<
h�P%pqB�.I<�d�̪�Q�D>)�D�/ʴ�{�ף�{��W���-�pXYVO��9T�����xl��p��q��1�g�E�r���u��c������}L� �!��|<v��q�"pEL�>0��H'�E��Ng@�%��w��(��tn�c>�zܦ�$5P��E�������Rq�� �w���W��6[S��iݎ-��1i7�3�ȱ��	!���45L�y�E���qY�O��)�^�(�f�*�6�[�X�;��W�ߵ�Q?�2Do=�����X�o��S"C!Fj������P�]
ڹV���i/Oew�<{��ߕ�X��cP�,_�-}W�h}l����6��@�wX�!�U9>�NC�w���#7M�[j�J�!"#�y�����o6?��w�2�,���Q��
��Q�I��ƚ~B��[�)�7����dp2ΔӢɏ�G+C(�SA�+�|���h3��A3�|�|��Tʒq�"
q�*K��k%/�����𤓪�o�`�]NXlxVHYEB    1853     810��U�N��,�vLC��@�Ph=��_��uyK�T�ݽz�G8�ߝa0<*����b(�Y@X8Ο�ѪGD�o|\]�4l�����Ҋ�������V)@�o�n�9�9�����;�c��qn�Zd|rgSNH�;.7nⵎd�� b��t�E�*�Q�+'P�Te)���C�X�Ǹ�����^j'�0��MP2u�[d}�4@(qP_��H�'���U:�ղ|�e�ș?�ZA��	ˡ�-�L�9@9���9�w���c���3���W��d&d�J�[��N�Q�����=���ѧٖxO�!��D���/��>�g�y��=e��'�Z�0:4m�x�
5�!��$l�>����������a��4%��9l����P�P~@�#~24��c�R��(��pBz�#,if��k �|"7�l?O�.����S4df5�P �z[7��:��f�N�(�������3Ϡ��đ����e,�zivI�Ӊ)��">�h���3
g��/���b��Z!�G5I����b.��.dwR�3������QMna��Hq��0�
j�^ܳ�9��癌2ȁ�r�1���w[ T��'�2��G�sx�Lt�ȭ�.������`�Nh���;݇��|7PI�P^�N�
۸uL)寎gn�h6�20�,�|����ϐ�K���H|衭B�Y��V���bm�2�JN��XPUM�$ԡ�x

���p���@!5f�^|.D�m����9�Do�a0�b�2�8��S�Y&�=�@�l(�S��.���B��Y{%>���ͮ�aUfE<�O־��y ��u��e��:���9�W��=.?���8dtT�u�9��k���x�ש�����RT�]���Ȯ #r�3B��ua�n�@�d��F�p*¯�l���י��*г���bh�5�!E�w���q��H2C�5I���z��A�@#^��5H�6f�caܨ�`�`p%���2�i�j��(����tr�s�8��;2�mT����#����~���Q��D�p�T���9<BS$E��M^A?V���V�7%�ޚ��x��'�R��A��B>��¨Zݡ�.B��i`^����͒�w��r>H������/�������o�!����?0Ư�jͥN����`��n��t��G�ki�#�O���״�M���ܖ(�XVT��'3�_�k��V.�imF>nj&��a*H,w���3���)��a=�Y}nˏ\�#���E��GQy�(�!��t`��b"e�{�O�i:��O���{o���}f���w`�kIW6:`rKEm��|�o�2,�Ê8 :\�kA:�*�yXQ<�z%-3:p�30�p-\;��<��� mOߍ�V(���P�v����3~��� ȠP��]��cĩ=�I�
�	���\U@9qA6�C	S����ף_��JB���M���$s�]�����<E`NBX���� ��u�^�Y���禠�9u��F�`��h��P�����q��7���~X���s'�1F|(���FR��RR���n���[\s�/�(�R���`.w�\��aR�
��q�����)MȲ�F~�3�X!=�sͲ�=$�#��K�\uB��Ǌ��@��pmVr�It rtl&�K��ȳ���Ԙ�d&V�>��Q#�M�S��r,�ZJ�?���v�-�8ph	f�upH
,�����}�صX6�]e����_�-ຏ�@'�4�4D���F�]�GS�� ������\҉=�J;/K���>Z8�g��b^� q��M�z��9�Z(���2�u=��"v�� ��ʶ[�k���sm�ZD�n�=p�M��wz��p5k�����3�s�U��AR2�G�~��YH��=rGyJ��@�ڍ�H�p����F��8�;�^�2�i���@b�u�!���2�DɎό��^�kA�h�F��/�:XZ���.͡P���&���N���k�E��~��{���Q����k	�7��B�(�"�