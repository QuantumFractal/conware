XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��qS��H�G�����K��#vu����CD�m����ҋ�N:�+��i����]C��$i�0`�kU�9���cX	�@݈)�{NH�!^N���k��~�nz�/��!��D�����L���86XM�� _�����K{�k5�3�{a�B��W��+�=�$=�ݾ�	{��L|��2X)j��7��Lm���ߵ���w�������s��^���׎&���7��u�m�����,(����A^96�if���1&B|���rEu�+�� Om,�z���\=:O��3�2��`Z�WF�������H�����UE���H%wFB�w3�z�r�#lO��:�R��fb�dj�����v~�Yc��yd���(q���\��K�9\I�_�Gc���C%a���������+Q����آ&Sb��L����n��C��g���l#�3��=I8S�)�~g;�N�KeJ�5����[+ى3���'���۱}}\Dx���S�HD�[C�M�����?���V
bznuYBbz֘���\�T�z�%�osj�CQ�gl46��>A���XHv�/� .|'��Q��fI�;���T%V�*��w�uJ6��P�/���*O�x.�
�^�I����˦}Es�1�\&���s��W��3�" Ҥ�=|������d:�Nis�HU�d�8_�8g�?d?aC7D+8�D���sI@��͚�Szi0"��8f+�=�ݔ[$E�i���Yq)��D���K4���y؄��?�F,uXlxVHYEB    6014    1840����K�kF�O���p��`_�O7;1g����!�]yA�vNd�!�4|����5�,�Zռ<p���� ��n�k˛��'T���>]* -K��i���<����%�Ҍy��;���A�j궭�l�\�Y)㠊�ALc�e��&0:��/�L��}A�r"��Ys�5%���&�#�9��pʷ��](���1?�9�e&[6 �[���{Eρ��LIV�J�R�7�ퟪf�Q/�o�/4�'cB2��h���V<%�ޞK
��������]v	���7��<o���CR�;~T/w&1Q'K.�i�Jo..&�/CQts:���^�QK�3�x�|z�X�ѻ���]#4�[��s�v�H���H���~���;o9I�x.�0e=Z^�w�m�-���nZ#�O��7�H��-7����4hd�e��N�.إ�7��dȌ�B���:L]���ڄJ"��)_�^���z��Z!r稻�(Ǣ��W�����%#H]�`#��vZ4�
�ǩ������j����Y>&��Fw, "�wk�Ǳ�J�I}_nNɁ����k|N~�.�د���S�1��	!�@Ǚ��\�ՙ[ˁi)7�]�Aj��������z	#�. �3��/ ��՘�:@y�c)^�2y�5�`�P.���m���g�O:Nzn��Z�����J.3-�5����e���ܥ��� #� X�<�`S3���fB���!�Z"��rc�������F�̞��pV��8z#tt�%r�뻾`yu��Y������ݛ�k��p��>��Lwi[�J�"��L�VR.7�V���1qM�|���K�꨻o9�"����&�M^k�:�n(2��cH��5�b0}	����i�&���ɶB\��w>+�G�}��_����O��].F���9��� b�a&�H92�[�-**"-��j/}�#�eh�x�i���߁B3�u%���;15��]��r����"\�� Ӿ0��bD��F�E;h�C�6]#��͗��TwcD:Cwo�M���}\�z�!���o��S��&Jw<5�31bv�M�)�Nx%���'�~�B#Pt[T�|�U��I�E�H?�u�����hU����M�"��+)��w�pd��x�P�� ���T��F(�~`�	�G Ad�d�	�A���b�2���Dɡ��X>�� ��U�ƽ�[��8?s�6�Q��YF�6�3y�1�t��H�>Z[�~���������GB��μ�	U���"+��9u3���)i��>�5��|+�2��ݨ��+&;P(�B3z�5L�~�c��q��*v>�����ymRѤ�&��p���'b��w3��b�P9wt�[��{���m�C/+���й��w�s��u��Ykx���xt&�uMTM�t�,Ճk��� �)�y�(s�_�4u]���1u*$�',�ʞ=K�f��hg��8{s�o�qR.�W�����pU�-���[�0��z$k�M�F[��c�b&���P��f(�L�74(;�	�u�����;��h�x+=���$D�ȹ��W3�3@S��O<�H� �~qlƥp�Ѹg��j��f0~Ɣ�"YǠ-:UH�yQ:�nO������v�=��%�t{ �����̌��8���>��*w\���7�R���`����X��������lЇN�$���-��Y$�ܾ���첪���0a���������6"pnX���Z�sn�g���mZ�|�9��%Q������(��K%���}xr�V�`�~TD]����ʳ���a�v�C�7ʫ5��J/%��I5\�H ,�8N��~";�Lc�$��w����l<,�^y�\V���_�E��c.�:�����FzkR��K-�#u;�[�	AP��<��m��`(Y��2� �2���ܴ�l&-�B�Ê�"�E��Q�A�	�y.V4�c"������M��c^~M�w���>F6Y� ۜC��jZ8�
С���$����É��ŃqYn>P�O�a���=� [)y�$!�z"��arY��k�Mkk=��
�iFy����+�t�f�7��岥g��
�[V(�	T�S<���2��:�kL �mH� �r1x4;_�W>>,�&5�`PP{��p��<~;���6M�g�]��)6Fx�1�b�S�	�pp
����_�N �6T�4�b53�0��VQj�|Be�[�䓯��rƆ�)��-�����J&t�Y+�~/��&��@H��&D�BjzD|��,��l@�H@8�O��o%}`���^G�^�%��DM�}��>4���0��ˆh:��E�	��� ��' �_F��aS�Zz� ��ͫ�m��.j�$��v��;��=w����O&>�yږ�ugQ>��Vj�i[)z�݀���(���}_Ә�K#YA�U�-�Li�_�YA�60�ơ�$��~|�,�����b@*$t���U+�~0OD0Z����2�ߣ	�hȘ���Je��R���7��S6U` U�����Acn<t~]�4��rCa�\E�DnG؋�R�j�"zڡo5u����a�M� ��PL�z��%{��,,��z��j�F�M��>"	A=����e�Ng|ܒ��$Ɲ��f�Ƶ��Ivd-����k�g�a#3�<�0�����.����N�	�M��5��F��#9�8�����B��������D���μ=���k��uDZ@�^~&����k�
��;t�Ž��~�)��Y�%��j�d�m��w8��p�����8�.e@�ߚ%�������W(�
:��}[�-\{����I�?�J0��6�ؾ�#]��`��FB1֪�iV�����.��+[�G���yS�Jܡ��K'�2NÝ�)��`}���S�9jT��y�m�xαz<�jnD�z�WN���t+:���M5S�`�*���oM�Zf���;,Xy����M�(C*��>��H���0�1��l#����tM8M��m fk����8�E��샏����L	��ٱ�/������,�> l��;���9�;�ɋZu���W�)�P�mg`��&�.���}��9E+ն��)�^�U?9]-�}7;�$h8�M1����~`SS�u�$雹�����Nl��,��u%Zf�%�|�ɦ����PB����ȅBKKv�� s*/��d	�r;�B�÷R�b%A�`d\��`%�������Y����+�<��x�n�Ş���V?'�{#��A3����2j6��d�:��q���PF^���!<Wa��br˽��xy��t��DP�7xt�V�� �!�5)gh�s�Q�qĠ+h��ue ��n����{*H�VЕ5�P�Ǡ�Ƒ�0ӎ#�\��K�2%�4���c���-���k|7��z���C�E|�,�V_7fL���V�N�8OۛA'��E.���Hh�v��7��2�~�L��=�XF�ΤV�na
�c��PM�)ъ�;��6H���|la��*s��K�U�8�WI!����r�20`k���S�8v"V�]�������?�2��>�^i�~������oUď�Z���M˳��!?"��F��Z�D�7$��S���CZ�_��t&�.���[�X?[F,��>�O��8�{��o1��
�- �m�m�H�+����EIz�G����i��K�w)������Ъ��&`�\�^����=:�Z�9S�CM]��5����2 ����mL���s2є�k�:S��Y>��2f�f��+�s��^��Z���g� p�#ɸ��kS�2�x��;��DD�;ʂ5�<�	J��>\Ҍj��X��3Y�@�B0#;֚��$�#5+���SR�����V����Z��Xy�RɯJ�͹�A�r 4l/l�b���6a(άG�aUtq�%��S<b<���]���9�g���hGgo��7m��Hx�!�<$&۩P���y��公�K�[aC��_�֯[pT֙�FyA�e��`�LZ�����n݂�	Q�)͝�c����a���^�@Ht!z�v>�X��F���
?�!o�rO��cy�*m��bí��K F�ڰ酆U<SnH>��9V��T!�b�����CX�;Y���w���aЬ��3�-S`l�-���-g*�_X�л��nօ�l��T+^����v�P8���z��w-`
��7�o��%0H	q8t5H̓C>��@���0x�Z)��ÒbW%�x���
9�&�aSOͿ<&/���K��2$-��)�J�Q ����w��m�jӉ�T�Z�b�
$�Ρ���>�&U!�$ �s5�W�-A9�՘�f��3
��t_��
�G�]�m䴒ݪ��P³P�)�/c�]Bu�۫rfe	S��v.Sx(�qu}����@&�o|����]g���h�ٍ�hB�e6q`Y6��z�E;��0䈍i�Rǃ���=�}e�^(�'Ϳ瀹��w����8�Y����<��w�ɿ"yX9lm�k^��5,Zz������H%?���6��̦JT�՚n7�}������Ni�ـ����3I�]����^��^#��]���O(��s>�j�1vH#��Vp�O�ӷ�"���|��˳�"0��蠲�"��=�(2��}�SQ�ܽ* X�jNZE�Մ�*�)�["��	��t�{A0[�;��C�`p.fN�ؐLU��Z>�b\�[@7�%Y+��23��:9�� �yH��Vpk���5�q��A,�]*����:H6���.{�l�7�����|�������2��X��q��i8�^�zkU(�ݡ����s�RifѰ��ԧβv)?igf��KJ=��Г�4��h��q$��a#:O�J���'��R�>U`�O�i+�\�����A`/�h7�Jee��������P$�?��V�C,B��a���8w��+�ք�P�vc�\\ �i�4�6�����0��Nw�QlqR0�	,�g1,Kd̖V�?��Ňz���ըO�k�=�x@N�嬦 �$	dnc��0	vb�"��Q	�W�|�5�W��2�P>���-���I��B�ް��M��GS���q�kAB�p�q�?"��mt��]�4,`���}�p���Ȍg�eZ���*�$��/4t�Z-��s�KD�1.��O��v��q���������R�g ���67�Cv=%T��c��S�q��0b�ڊJ�����+.���<~1Mڑш�[�Z������9$��K����7!v��,p���5�m�fR��t`��Q�(�n�y[��{�t�
B�Ղ�N?M���K�{j�������y��$��𺾪���j�y�ȷ�ۍ����̻Y�^L�"�z�b����`k����}&)��#��y���+���t1+���[�c�Pr�^G�ļm���	�������X'��cj`.�9�{�:�1'ղÞ8�9��S0��.�O_	s/AA���EG��̑+:3�N�{
ͭ|�Ss����EUε�R_-��n�Ş�@~��_$��Ƨ��H�͇)��e�ut�E�T��g�Y�(s$��5D7��D/u��K5��SM�홸༄����l�i]��?2�w���UhŘ�-W��j��sm����)�l�޹�h��+qK�Ѿ]?�ĸɃO[L*�6�4t|w�gr���	,-�.��+|I�D�U�f�Ã9D�}.`p�S[9��Xs1���4��	��RRWl�
�;��+j�]ƌM���>��0�=�����F�0�H��|֧\涑(_����*����6(�\�]��ZL;ޤR�	������/�} /ʏ��;&T���&��W�ܢ�����i��fI��вK����s�),�d:*L|����/�DX�1{/�Z;c� ��u�H�e{�,���0J�Ӡ�+�tl�;�,g����,M��7#��,ܰ�2����p��L(�Q��\/�B+|=�WTՊb����S ������١h�[2'ҟ��u�ٴ\{?�΃a��D׷�">)�7��+�<[�u�%�B�d�S:���߽;��R8������4���V�����2"�Ss����lP3.��[sԆNVq6����rd���������1�Ī�����Pƅ�����t|z��%�@��� ̆M