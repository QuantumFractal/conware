XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���xi�BYC��O8�V�^n��
��6jXs-���/��h���q8jU[�%XL?Y�R��@iT(�
P�(�v>�sn���o�Ë��$�(�F��MW��}ʤ��]­ȋp(���z��q2�u~q�+��OR5Z�=َ��������<�j�@R]T�i���,��O�^ߵX�x6!�_��Wl_�ĉkhNv�:K��Tf4@[|UĴ�ЫD�c����!l���2v���8X�
b�J��S�cX�`�W@%��0�i����.R塛�."�Ӡ_���-}��C#�"v"�����Mb`;�O~�eEܭB�hi!���g4��ؘ.s^��\Q>+���F.��鎽��h�So+s�:�Fb�t"��h�"�����͸�1m�ִ[9�Ђ&�H��ڇ���r35v���F)h�S܆%�+�&z� ʤ�5�3-��Ȉ�ݕ��dH�6{�N��/����i��߲�${\c�C6�QΛ9��LE�㊟K��R��ЮP�'I���^�d��ׯ��p�`J��l5��Ǉ�CJ�20��8����C��.h�w<?�[=��w�$��&ocS�ĸ�m�$!�مt�D��t�V��H����y9G�5M��l���S	N-�%t*G�}���t�q��Mx7��v^�pꕋ�9�=v�N3��13-��&�P�"�C�疉����o �t@i�����-�D~d$���k� Jsa���	�=t�Õ�oG�T{q�gY��Pd0f����&�\�^s��<x�5�XlxVHYEB    6346    1790_�#������_���<b�����6|&;��������D}�C��-D��"|�e�r$p�h6ۏ.�fz�@i�a�L�,�[�>@f�*ۭ�᝴X	�bzL*qI}:�/B_�b,�5�7�c�5x[l���LEj�,�IT�5G�.k�H������&,�>����;K��a7�<�8i"�ҧCB�5jzc�t��(��k���f��eT5n����fm��nی/2��Ѧ�FÃ�Ʊk��W�cݔj�H��9�J��xΑI�� 7�/�p�����s�6 
L�UD8�D�>�l�֋���N�P8�>{��EO�z3�8d];Dho�d�2��T���&#!�I�9q�ڭ13a�E?ZS����9#5�>u�.�8v�=:y3�U+z�0xSN�L����]~ޛi��=���;�(\1t�p��oA}N��FC[�Ԉ��Ό9��r�5�t���Vg��Q��[�`Q#y�X=d�ۅ*�;�+ ��:C���� �FMB;�6�=Tӯ�����ˑ��3<��_g9Y��Xx�X@6��l�\�џ�C&�E���L�R׮���l��ۻM,
<����H4
�ycL�$0�|�T0���[��az��{t�Z��f��K~6�֠�_�V(?B�I��`�Y��yȱd��ܞp�-I�͎)�M���gS��e�M`UȖ5o¶	U�e���f#K����
䫓�u�}�^���g�������Z�
*�����-^փ�{���8���>ViJ2k� �4>b�e�����u%�����S��
����������i����|�Q���+O��hb�X޴�����({-�c��z9�q[��#RR��������@uV�ma��P�v��ŏ>l��wA��̹�*��Q��:��J@��5�SǮ���ϴ��+E�y~��a�o54��NMO=�f1W�4���W��9�����\�;�cܖ�g��g���O��[�Nqƀ�U���d苎VWx:����&#3�ȖB|�:Eg7��;Ү4!��ޱ/,�����j�l��'�
�w݌@�<�f@}'�����pR��OΪ�C�.u<Z w6��q�����wB^�"������VD�g?+��6�}�EZ�L���+?��?1l6���4L��
�
�d��_����xe &��m�lm�]�QW�LLHQ�J���&�F@!�bp�9S��~�3P^�_����O`}x<Z��lc)���ڼ-�2=�V���e[��΍���:�����4r��I�[>�\�Ix�nb�����%>`���<kh�;����M�؅k�ȒoC��kn��$�r$���O�^YE��/�l!��s���Z��7��ԠZ��g�?����)�%`R<�.H�)���n��=����x99"�y)&��ڙ����ܿ$w5f5/�q�	�����D6�h���`�t�R�t�;KU�$Έ��+���Yț!��m�I"t�6CU���<o�h�X9�P�9j]��
/!: 4�do>�f�D�&H�V�6�l��[���2�1,�Uu�O��|�S����� ���D�m��b<�C�>�!��
�{���`��0���f"�n+� ��>�W�ҳ����*� q����ʪ����] �/�î��Y��E?Y��~Ƚ$�qһ����-Z�iuTP4/7ޑ�qJ�|,ßFrsg��	��_��I�����`�[�����2��d��>Fܖn|T;G�7�
�W	=eKq�DkU���2m9q�H��Kz�}�����x�#�ںk�6n�����~W��|�s��ǃ���] z�L��g
��q���w㽪�� p4V"��}_]�*}^XJ@/�.�$d��<���#Ԙ��	��0NW��2�����`v��v}YAFmэ��Bn]YTG�oMN�Y�@����16ƾ��)�x�:�����FWꘝH�v��,m���B3_j���(�3��"��<끇�&:h5�C)�"%��M4����#@2YvJ��J.׵$4�"X*q��f2��q!�wOyP�D2Z慟D,��<r�>.��h�����p4�n��s^0��V͖vY�gm�99eS+g�/������j<� ���V�;Xꦱ�#��?�}u��ә��ah����=�c���v�[��OP�d���L�V��ҧ�+@%j,��n���7H��@�/dwF8�O�̈`x�odh����D��@�L�L����"� /cٞq}�ߍ=�>�ß��iq�YߗDo��z�e�zq�xArE弱+�qH�[:Ϸ ��;b�we�1'{�V�M�:�%��������^v�El�%��#M����
\�������˧>��5���X�<�F��C���ފ� �Me��{�]k��E|����?kّ�$�ӛ��4��}q�!N��[����b�~n��,�5Y5�[o��W�j����M,n~�ڎ�7o��F�_%g|��)��N�Kv1>�� ޒ'��!mM�h���u�B�*1Y�Qs�Jr��)�]HFd���ї������^_���Ҍ&o��=��8�9�D�w���:��eV���Ub0 .��ǖ�.��/�` �G2�KU`}�$0��r
>ww���>$o�2�wR��_�@�`� �~5���-�V�� �i�	��6G�cE7ú��fj�-��I�BaA�g�"�"�x���$:gI��
wjX�X�^�1�j̍��X��	�T	v�s�AGj���R��0C�a*+L�=�w/y�<���i[�{P��p�W=Y�[�5��Ts7�}�ynR��
�5��5�Sĵ?��6�>_dȉ �����w����	���I�5�<�eRӯ���c ����B����0u��fQS�7�0!�g}4Ѧ��	�Z�:p�E�К�Z�q-:�%yh�`5�M�\^@���㷭�Ʃ�s^R�lɌ�f#��Μ�\�ö�y�r3�7�.%���+�&�VZ �<�
�t���q�B~���d���1n������p+���%�hb<@���P\�ҵj�%���L.����}rܥ1ݘx��3��e��3d|�1�p��Rl����e]�~��K�|un��UU�c�@| ~"@�!��ei=q)���MY~5R�u��I|W>1�)[��Zm�������8-; `�U$����w�l�NT/6\�q�t�f�	��G�`�%�� ���m��N��E�n@> ��M��pV.m��D�O|3;���UZ���s(�U��g�۸����)X�Y�7+�� �S���J
6 s6_��m��y\tO�\��({�l��b��u�{E�2'�6�.����?`.��R�A�z%��	��Q�(�܈B��hD殍��|L��5R���Ư%vIF�������5i��h��8j~�ku%fE��W���Vr�T=mFɆ��6lu+�^��=ˆ��`�]��N'��ڸs�j�]։|J�J��h�o�GSm��X zm�1��0Z�)���6ss�6���m��J׳>��Q�68��n�w�X7�ϟ�͉u@�����,��D*i]�)��S�_:�:o�rӢ���0dC�q։Ԑԕ�4�yl
��;��4iv�������/M�PC ַ��$��(r̶�d�))h_��l�A|g#x����^>@4KVB���̃�����ΧI8�w��R'�m���y�G��h�Ѻ�ےx�9/�v?o7�<��v��,��"�_�8Sp)D�Po�l���
#K��jP7� &���*T`�=��ir/���z&� ���l��Z҃nn�R>p]l��׾�N�%u����0��t�b�[�Zef�٘i$mw�Y�K���ܑ;V�r"mS㞆�%uI���Wq���J1���"*N]h�FeN��x�U��k�΋o4�i�2�~$��7uԱ1�{��@|>�A�wؠ��$m��u���pu�9d�����?�~��[D3�����鬈�#S�urd�>m;��in����֜�:G`I��f+^D�<��0`=)�2턏�t� �sk	����e��y��ED�������d�:K�(:�%e��+n3VO��LY/��Q��Iᴄ���^^��\66��L�w�l��(�]�f�Ù���i�l��f��A~�.����*�����ѱG��/46��6��uf�~qȐNo���������lW��[�$�L��'
@��B㷞|�WFVᖧ)�-hi�ʆ������x�]J���tW�u��bJTX�R����\f*�V�x�l��/-(Z���$0�(��;�-�$XAK�।�@�L���$���}`\��H��m�&}�度� �*9Tu�QE$c���P7k��0
I��<,�)e��"��3�Ύ`�?͂ҭ�#�)S$�������x쀝�'���~^V�^$-m�H��a�[\���)���2 "����y��ԝ4h�Ղ�W$��
�R?�5va�����P\�����<�ҏ�f���ZNC��'v,ty��:H��r8�1ġ�M�sT+��'Nǽ�8�n�/=��Jb���o��lA뢐�s���7��峠3�~n�K0u��+�f�'�$�NC��H$�#�f�w�lgE/u~�l`��b\���1�M%��+��`{J�R".����'����a�����ݝ���#�K�!j6��G�C�l%1�mD\wM��s �Mi���ʛ��G�A4}s����,��O:���Π��]F���>fJ��:`��>ӨewK=��U:�gG�����Z�P��Uc�s��T\A����G[�qy��VQ�����3��I'��a�����}�'���;z8�s�&d�o�nY�Dz�v��G�W�.�_n�q�I!�@�C*o79
X�#`��>ц0l�Cy��	��
��?�E�e9VG�����[���ϳ��J�㙐����X���>7���J��X	�va����m DgG,�fS���	_�"��oCss���v�Z�W����$]���S֜�=��`�F��LL���P瓕��Ʌro�������X>Θ���cWxI��w�e!���k����ݧ������-z�j���L���4Xm�n��ic�ȃ�` E>�\���s~-*�ب6���?D�q�%m�=�<aЀQ��p���M�h�{^�	L�yx�!�����}k8�GG(��������#�^RxCD+%j|l��~վ�]�����~-`AW���g�4 ��o��,�*�-k1��(��V1{�����g�~9��7��?=��3��%�,�@%�N�'��OG�%`>k#�:���c0�w�����ù�"uUO�)Ru1����Y0��V�\:���ɞ��:�`#@�����8[�2,��qV(NC�2�W�nP���ܵvE�
̓���-W�8Q��r`��~m6�	���(ɥ�l�Ȉ�q��0b�w���'a������$�PGan �9�5Z R���mC��L���r�{��	��h��UWez��Oɵ��
�|r��L����qF\dl����$�/Θ��L�>$�|�����
��b/�oT���Qi�5�J+���Ш�{=��Bh�]�Ȋ��$��M9m�M0䦪��²���e��A��1؀�۵!�^�T���s�\�{0��^�W����qڭ�M������t���e�W�DhY��:~�����G5��%yV��p������-�:?W�����u�
�r?W���v*�����w��K��(XR�2��Vr�s�ul����s(�|tO�x ��^��j��Ǜ3�ũ��Eع��.vɲ�p+5����`'~E�sĎ�3��������o���h�T��\����⣻�.c���Waה� #y�DO���:��P�H謥`��{���/����T�ŴӴ�{��+�t	�����J��F;�[�b���	�aT�/����|\Ωa<[gHb��2e��t�L�