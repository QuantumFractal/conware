XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���r*EO�_P5�6�Շ$z�*2������p.yMQ���n=�FCP���[�vX�⋑�`f��p0��9������'M�BS��	~��o%<p����(��e���P���fm�e�F��ܤ�M蹙���iʱ��pٝp ��ܔ��F�ZQ;iFd��C���h�����Ձ��׎έ��}/G�XY'Ԧ	���6��s+;~�g�_1�ˠ5��g�>�h�cs��Y`V�S��;�c(��̛�Z�ۻ!�����ޕ�*t�6bb�.iq�t�=��A-�����J>	�P��C"m��Q+�� �vOW�(Ig��J0�֊7��s��&�%� L�'��Tຂ����o���0 ��s��b:<�/���xz�_��'<Ń��>L����$ǝ�Uq��>�c1���@��X�!aøH�	C��łh��Y x�Ζ�K#�}33��� #��UM+�8�nj��߼J)g�j�IЂ��<������y �O?�}M"�e�&sa#U�d��کd;W"���)������8���|�����^����P�vjOm�]�W�r5���S^x5��x�_���\�(�d��@�':	�ǎ�]��E�	���7F���y{]��	�S�^�X�;�lۗ�*��4�xDP��&5�,1���N$��Dŗ���W�����x_��;��q�ݙ�:SOf�<�����O��GR	c~beĀ+�V�k|G���Y�D���%-�B�]��6���e������~M����XlxVHYEB    95d3    18d0��˗;٠%��o�;2�]�#?���	c��㥎u��y�:�];���p�TJ$�n������P� [BOΦ� ����k�0�sIug��23��<u�Rׇ�}+��/�U�I���'Q,ڪ���k��!l�Wݰ9\0ݺ��ڛ��V���k;5��l�����i�����K�]���\�\�"��#,�E�̓r{Q�cKr�0�ׯ�F���qe��<�Fٶ�L�k�q5oH�'��&���E�\7�O��2�\�{�/V�-�h$؂�7L�AN��䜳f���܊�2��$*͡�+���c[z��g�t�\�c�$�Z���B�/Zl���ZSW���M�o����B�y{%���?g��Q�nQ�@�eG�����N3�y��uĳ�����C�~h��� <�;�*	���Rc���Wp��p�شV_RH�X�OH#�oX��ᇃ1�sv�^�Y"<$�	����9<H�Dc�*��]��;B�Eᤖ�/������9���ȇ2�
�%?�ۓm�_���lԡ�U����ʌ��;0����˕䫴�Q�w$i����Q`�3.�ХPk~oA�(o��򒌂U�O����vs�3)o�TK:�Ol�l��<E&@~��$ǑB��&�I�PR���/V�-�����Qq D�O�i��ݹf����$�Y�{œ�^����ЙYV�3o.3�"�$Ng	�x����������	O�R�Zi����}��Y8e*�^B�2޼��D��J��������;��\�>*�b�V�(4A��g��-����I*3���>[)c}JP���L��Tߢ �p¶gG/�o�x8p���Ŝ��<���X�jh�M%^�{��f�dvv�
��F��!���t!a�f�]
���FM��y'��ο��g�k�f��a/������˦6�W8��xKWRVX&%�gre��ys����������{�~8��}{G�M�Z��ѦLX/���j+J��:��K�y�86R��EZ9]V�8.D�rHS�=Dč_[����B�� �=~����Z�m6�CH
�����H�ۆm��,�\H�pA
ayU{g�	k����L��(�O�I�`A!�'$�_�]t4�5��������"�+��qJGS*�}K�_�.CE&^l�ݝ]WؠD�V�5������,IՒ�� ��]��!�0�_�2>d�_���8L��V}Z�S����� r�d��2?܃3����٘�Ub��Nژ�π�0',(�����}�R��Z��H�2�n�O	��id�#QK+��r"Qj�z��v���1��WTȬ悉ΰ�JߋɦYԘ�k���?s��o��h�CV�cH��?tn��[l�������~�D�[<.|3!H����P����[��ۏe6ߴ��\Ӽ��9��m�'b��.��ǉ����˷�NB�ڕ��x�y�@�/�v��y)�xц�&?"�K����w��љ�޶�t[�7�{��
�J�A�.쭋�OX�A��ˑ����I8�Kl<D�&�!�����i��,>�
�c{��HV������1���s����<�Tz;�)�1[(��~Q��
��#�H���K��FK�$�@z���O�NƠ
�^�Ж�;�:!��#B�Ra�mf��׻V��Y���ݧ�|��	c��W�Jt��4�5V�_@�#��t�)�4��{��+�XF7ծ0�w�f���
�{��1��#�
4w� �V��{��v�9��dɒ/WbM;#�szI���z��ŪU팁Ӧy������ ��2����b�B���&}��7U���k�P����@����N�$��5@h{0����
�"l�S�%x:�r���88ۙ[+�Zzq�^W���	�����D�|�4&���gN�U�p�k��]��-�EQ��U�3��Rȱ#�y�� $k0݅�L��и�aZ4�=C�8�4Ѽqwb(�o�L�� ����~k�d�;�{|r�����<�2�.���q�m�u�8ƕD�=P��6^���2t
w%�Ė?��Bhc�O���KiLW�&�}6$r���lU��k������;oŝj�v~*ti8yžL7�JA��cwx ���A{:����k`e՜i�^�I@�.]����]����46������0�8ΕV�<e@����Kk'Ҫs٥-'Nq�
x�}���K���vt<Xh���*��d6�/Y����;��'m���$��+�~�d@)�;�ꩌk'r��^�Y8�fwp^\	W��?i#�@�|(Ej춠u��{>��$�;�1Y��!����=���.��}�{i��|͖V�Ζ'�#r���<��6ϰ�R���FH&P]<GpDG"��X��#�NQ��E.y�uW�kT#یd��蟔��(�����H:H���l�0.� ����Q��rT�-�s���,�p�hU[�٣�5�U~�x�%���;@Kс��Ќ#��ǺG`N���/�!$�r���~ �A��ӟ{ΉL���t06@��v��d(�4�u���W�I��p��*�cy��P�r�	H��dsJ@z7��h���{f��}�� ���l�+bZbaQ���a�\O����j3��S~�B����p�9�1�j�ۨ�z�r���&I	?��4�c�h�R3O�R)~����0U��$
s�7��?��c�*���OA�ڿjիm���3�Gԗ>���af�5][M�f�6�fo�(2���=-��x�G7�"����I
Tu�a%D�w�r; �k�rhv�*�K
oy���Q�q�xS�:�۸�D��,Sݬf�*'�5�.߀�"�=���̅��h(�/O�|`����\u;3ۧ�>��Z۞�aNw?�)��\��^�7���u5o`�s�ڬ]]�9J������jX �X6[$E0�c1��1�o@�U<-m����^�/�.��B�:ł�^j�d`y����w�G��t	��˖�qW����ő��ݍ$-�Y�zB��S:���,V,�7�M�� ����>���,{����+ب����J��xU�	ў�,ۑ7�- �Y��2pVE!���DH����%X�"��ݗV��:�aZq,.ǐN�3G�����C Ѽv�EF&TI"]�Č?���j�����z�yl�HR�B |�`}F�W����W�P_a�yCPr=�H���Y�ڡ�w0�3�:�zd���޻�mu��H�r��˛M� �q�؅��ƙ(j��j�>�+;*�̓T��S�x�]:������ԡ����j]��Cee��ƃ�߿r����m/�e�WV��������b�7�2�Sn�ץĞ��ѡ���#y���aK:�\��s9��#�14IRc��+�W=�e�x��+=B-�G��#��	�v|A�t3�E�g���}�Pw�?�.�f�Gǐ�M�(A域 m!�Ҁ��B ��<LST�evA�x��@�Z��S��&����
� ɍR8��] �tbpHQ�q����4dz��.�Y ,k� s���,@��2��W�&-� ���}�����//3~%xE���R��@�zZɛF��k��!��	Sp��>N�NMH�����<.�N��q.���, "]��B��������y�e�R[�Tޘplv��Q�a��R�]>
7p�U=H��S��#3���<�A"�� T����h�F�r���*�	 a���S�* ��oPŕ3��%!:yϸM[6�b��F�!���9V�q0���~׽��p���*"Y��8oMR�I�6>��1�ŋ��!=�w�3�Ν��ƕs�*���t���hH~L�����Xxe>̷Wm��E."8@�ˉX�n�e�N��lq�h+Ox�����_s+=4ߏ�2����U~��X�����b�eg��V���G��]���r�'�0/��ABʳcoٍ#&㼬06�pz7��]�&��ܫ]�A_��T�k�E-�f*��k�� ���O�r	P9A���#�
�_c(�;����4���:��U�����H��ڽ�� ��Ů]�-,l<��7&Λ�0�Ӊ4И��`��[�L�"���N+�GQ����h��3�yk\�iq���6�V���3��%omt4VD@�L�ޠ������-��]��<�ɝ8�%�T'V!�Z��C�^���@9�h��F@�1��m`i�,>�Tj�? V�C�P)��eL��:�C�:�Ug��}6.�ﴀv��a|�;��t�j^��G� r�|Q���ɣp��~�h�_����X%�@6�PZ2�67S��OK���X85,�G�LoQ�{�v���-3.���`���!�W�Q� D��g�Y���[	���¼���؄q��O�zG4��M#���g>W:�
)�( W��$f1�Zj���Ԛ�;��vL�/���d+��\iA$����~���"����-��)��*uT�v�@�<.�ǉ�\����E��v����ڢe�ELR�>����������?���G[����
Sa�g3�BCD~�'8� �
5r��.���a�g�M)�&�"#��Ń���"aJy?5P����mh�ORHq��ߵ���-��������/V_ |�2E%�%�E�a��(��DE��y)�ڢ��/�1�	��&�F6/$Q8�d�Ci\��jWA\�=*kw,I������3�YH�2��*)�p_��\SP��B�.���K�I^`���Ϊ�V�-�̖�pQѝ	���d����|�|�W�0���b4�
����gno�i�����A�o��=������/45�o�;t�TwՋq2�u7LQ;�I�ML��ą��-2kQ��W���t*�	�Blќ|"Z#}�� �����i�5n�k?�����fUcJ u���BJAV�E�dt��+Ɣ���B��?K!����{���	���8��{,0߸Ȏ�C�LJd�4���Z��F� ���ϝ�p��qQ��\a�?i��.x�J�_����� �H�r���P�5OĨw�QOC����U�ȝ{�~��Mx(GS��1�a�B�Gm�!���#mr ,�����!��	:��J�f�j���(��QR�~�NxRVu�I��,o��k)�
=��V^LS�r��-ovPS{�nWhRY�����(��R���҈Ь=^3���C*�@M��T|W��P�UlH���7��8X}��<-���m�p}�{|�z'�M/s�v/�}����D���P��!�W�ȍGܚ� Ü���X|������A�V���{����Ct���"G�n����p��E:\.���s�e�{�!)����Q����f��I�g�Pp�U�B�9�{�^Qp���1��&z疇�0��Q��/P>�ߏ
g>���1ذ >nb��*���������ce�@s�5�95���O��j�ޟ���h�����	���77v��	� �^�ǲ;͛;�A%�r�	��z��E^RY��y<����@��ϵ3��$e/�`�~b_M��{T��}^5Rmn�'pؔ)�l`k�X�_S�����7��tkz��^4%b)�u�I��9�"\_��l]�A����_H�NU� uh�
�C�W���UN����q�/�\��%5ٶԂ��p���ʫ���S��lk���[{�e��gn%�S��_R\�T�? hW+b��ky'eu����'p+����	U`���n�JqD����Î�u��֤r 9
>��2���j��ݥ;��!@�����F���1�~CB���	��Hܤ�.HN���Do/�-2���"� �m�ID7`��<O���!�!��qTڙ�\����>���N����S����������)z��^�O�7��پ�:v_�E��2��/,
�n��Mq����v K��پ�cң2 ˸|���T������T�K>^}X]Z�^S�;-k��CoN�a�.��R��k��S;	)�;b3�6�=GH%#,
��Y��m���t7�q���ý�$n~�����4�$!�d��"�G���dgX����U��W��b�MµXݼ�B�ؔH؋4�z:�a��=[�Lϒ�d�̚�J�"9��vLa��:v���ݕ���(d��S�[4aS7��^n`e���%���#B�4Ȣ���V�Ro�Hɫ[�S�5� A�������H��p���q`oz��G���q�<�G�.��N��)�p��-��`���'����G�a'��ιWu��~0͖X�4$wDag$�k�vI�h�A��9���S�|,��0p4��gy��0��q�����S���F�������ǐ���d5os�K�>pY;
���0W��g�