XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���,c�b0���UQ���jS��̅�1�dU��N�[�� ��~o�4�1�(��V�q��o����T� ��z�]�Y$GΪ�9SFv�����|⽯C����t��2�� �`�(!�=�S�;��Д���X��E��Qݹ�H�8K�~��[#�sa9�c�� PjMǾӛI.���&�t�)T}�,�����I���ϏAڋ��v`Ƃ`"6�l���>�� �/� f4X�X2*S����Ĭ��D:?A�����o�GG�g/�hy��⪛�	E�K
:GX>�Y�* ���h}f��Bm,x��-	
�������Z���J�͙���F_�r�D|bi� ���y��_!�G�z��Z�}��Wy)���s��?�w��r��5(F���d��U�|o�X.��gF$@{e��&�0�ٕ�1�@�lr��L��W*��d�)��nd:�i
��s��*8(��W:�(�`,>�,�ު������K���̨��C�n�P��Gq�3��!��e�����P�Q���R�lC�i1x��v�ZI�^
��WO����{h;�c��S�N�}�͔R~E��
N�iG

t42�XL��'mfD����rK%tFW��m��F�n�'Z�g��y6�0�6%�4QMT7��@��0�*��UF��J��3ᚅQd�d��=�-r���\,��`�>Lj*K��m�W%�$��m5<�^= q�l�蹐r,�a��_!v���$��c�-/Q"XlxVHYEB    fa00    2040��8��FG�\����?->�/�P-�A\x~�O�zb�ܝ�<һkb�h�O>Pv�g	�?�Zv&�YK&_�.�z����J�Q;��/�`��ٍK��4Ky$MTeI�.%�zș�f�k��'W>�����;� 91�Ĵ�́�Pq�U��;��̧
�*G�H]�@�?�i��C����B#��;5H��ޫ�m�$<$I��$I~7��A�m��ɍx���}}������&N(�� ��b��������ԗl�y>@M���\����9�eY��*�!XQ�[��"/��܅�����a7IB��@��8��Kl�˳lR͢)x���B����M�~hp�S�)s`}"9��@D����~�L��CQXѻ#������@�Ӷ݇���f���D� ^!�3!"e�+:C�?D�_JGjJ��r�N�Wn�𸐟���Tp>	�ծL(�:���U�M(�ngy�/��^�d����,/h���;H�X_���c�]��E��� �6��L�i�u�E���s@D���윋򳯬/�	���7�irj��� �5f�]W�(�m��v~.N��J;����R��筰7vzlИ��I�{�CJ�Eo�ya�o�D����i�Nž�fT���I�B�_g_��ˈ��_�-ƉRa��]ʋ2���0�lO�b�(�p�v���U\(WA7��}н(���	���@��,���n$c9��C�(�a]�^�;L��="M1���r�0��$�+��P:GV�RQ�CjQ��`�h�Z���*}���p-�O��E�P�-"�siN��z��WI(�_�.� ��^:UL�Y]��D�r
���E�+�7X2�D�&�z��$����b�O���|�C|�{rr�)�a�L�\ZOJ��#�Y�v�MѬq�2���:�wQ�aGٲ�����N�@�!�Ȓ��,���(�R#W	UQ�Ŀ�J�q]���".#�|_D��-YV������x|���$�ގ�!��I�ͱ!�؇�'�ʹm�yi�5�s������ME��B�I��1a��cIr���cm[{��Jt���l�yiq�����m,��v�e�~����z&<*Ps��7)�ƙC휊�2�<:έ��i�?�(Kev�ۚ�k�T�������1�?`2����~Q��Z����G��X�PoA�� ))܏�n=ߍ��+�ߤ�0j�60\�U�U��k���I��N����O�e�������{�6��*d'���-P�KS�-_�����z#g���U�&xD��/0�wTgy	e��ļBg;�2H��:�w᥀�7O,"kv���-��˒r9�g�_�Z�P�U֔�O��-?<}�7��KE�}�r+,<h7���<"q�[zI��hz�r��)�������\d��]q&�-��~���5��TK�gĉ(g��{u1'\*a*�������b�W��|�l�����}�ҕ�9�1ȒJo��V�IP��i)�G��*�t�DIsK�wdF��0���	ɥ��k�!|^�֐i�≀4>�fCܯ�@�����I�z����	���k��R��h���,;�D�Eƍ�)xH�O-;��qIHN�q��kȺ&m���e�qz�r.�J��LJ�q���--��I��pK��I\�L-�1e����L���e*Q.�>r��N���%b�R?!z�a��y��?b�n �Fc��1Lk2\g4��+������HV����G'=�&wO|ȉ9����Q���s=�A��(���V��iӉsj����\ą�ޝ����X�B+���/�����b$������Y�V�W?�|}�WUɏ�˜A;C���y3���kp���ņI�'y���oW*둗v^-�@�B���sH�X'w3�[�<Ki<=��8k���u6��{�Ee�Q�WB�b�b��BU��s[Q�d�x���Q/iO�o-�r�;k3�Xا=.�Z���`L4uJc���cME�����^��mhМ�/��8�C�7*%s�����*��Z�I;�&r� ���a\@�+��A�)�j��~��%��C�A;΋\�����Ƅ]x�Icu���+BR� �Y�K���OnѦ}�ƪ�H�0�/ɏ&*ű��H�v��K�8�::�ٓ�H����|y@�kR�YW����)*��������y �uJ�Hf�6e�I^��9������+��H��.�vC�̞VP��vz�C��� r]��8< ��G��~���� �ϔ��&b�G;��&�݊���h���8��Mʦ@�����!��}q��"w
��S��i�eﳃqڱ�>�����ǡ���L��>#o'�|�8���άK��S�b��@��VUB7�'C�e��[=���;'Ƚ��Q���Ա��L?���~в|��<�ѩ�M�"�F7��s��t����	l��0蟖9���T�Y������OU�u/�T�7�3=nW��x���p����R���K6�J�Y�'o�(x)��^T�

t1�pA�$���y-23���o�{LY2�<��%R_��љS�t��T[$6�`B�H�L��B�����L��i�y˶7�8[~Ŀ�o3�Fx)l���e\��:Ļ,^:�� �l|C�
5���+S���I����?���?�T�.BՄ�;�m�>�GKR�G;��t�*�,Yz�ʴǢ� �>L�����ʹ뒓 _��� �ٕ��0U`�[xh�Sɐ�hlͻ�\k5GO$�Y�Ļ&��T���-An����>Y����,k�G�І�����G�	r&-�Ȝ2k@َ���� ݏ�g�G��I�bM�Zٴ9J���?h��պ��sxCˣ���O?${���e�����Q��xI�ÿ� �fǋ<S�������B�SF�=��~��R�+�%��n/��b	Cd�"�a�3��bhWۄ�[�2�s�W���]��&d��:��H C ¯aN��Rc�m�k֧�sq�c���M�,|'�YN��v �}@CZ �lTI�G+|_	R0�ס��d>a��*v�
M�(zm؞^F=0��h�C��-F���8����B��T�?z�����S+?���N1Q:Ra�������M>�����N�(�/��r��ݽ�K���������ȶL�)��b�qPU��Ep�_	���ҷy��3�Ǵ�	/KL������]L���w=�|ᭈ+� �ɷ�#ʵ�`i�� и��g�D������1c.��J��ze�}!j ������߮eȠ�qg�b�V�X�b���w��em�:B7Z}�J��U7�� $&�#?>��;5���L�^�����k�u�n�Z�	�\�Z$j��_|Y���J{�+�\S���J��h<��N�O|�%��U�'ʅoO�8��j�0 �7#|�"�j51���>_xN���#<�gj��6�<"��G�*��Y�&h���5>�U5T���ҥ~�N���_1���>La�Iwu�u ���r kK��\ �,ƻ1���'����F�I�����oR���_zk,�UHbJc�ܭQ��U�w!�M��M1?�v�m��?\����2���7ܶ����^!�C�qr{�����Lp�`������f̴�$<T�.�j�{d��f�;@A#mҮ��ɠy^�l�S�ܝb�yq�	��qK���}}B�<������L3��&�ߪmrÒj�f��٘����u��q�0|ubd�>�h�Y��R� ~R�UC�$U2BR���7�?t�3Gn����0�_���h�~�Hv�ƅa�˱�����|HZ+6},��7������Xǀ}@�`0'_ѧ���+���>Tr�	�}�6.���&�>K�A�QkO~����L'���2�����C�^��w�2��(e����mϐ��!��V��[�������'�z�`�*�|Wi;�Y8�+ n��S�)�3!ѩ�风�A��K��R����ŧ�X�����HP�H9l�]}5dw�l�ݳ� ����r�ٜ_6���R2a����[`�;cA�#�M�Q���8�=�����1�8@|`��o�$C����=,����{k��[���:C�!����CN�)���v3Q�w����c ��{�SشS��^�����/����~ ���$�K���߄wP���`f�I�����F���hY�P2k{�*M0AC��E��`�'�q��9�y�Mׄ������;��Y��pj~(k�I����"5�\dg B&���I�d��PuYJ�rqDܠ¶��~r�{��rE;�P�����KO�cM�]���U�'��1C�&dq������v��Y��'%��?�ˌ��j�@�U�U$�V=�)�ӧ�6�g�I�]Bt��*�4qU�T��he'#��݋ɕ���<c�.Qji?Ɏڑv���1�?8��DZ|5��@r��h#櫙0d�,9!�(_Fy�(2�{�fFi;e~�	�F{���s�S&oUT3�V�޹I��C邏���6�נX�Im�h�M�1WG�)��uOSkݰ����6���}Y�O�+������Zz�dE��*� ��q�=1�&�2 QRW����Oz�&h���M]��z_V���>2�Y=bo!b�mh蘏��k�$<�#Y���?(�f��%����� �(#KPΈ�H_Ly�ݍ��$��|c�y�_d��t��Z��-�}�����
�I�&>`H���-��}iH���r2��V
^_�{|Z8�2څx�ۥ��,�CJ`�X��H4�y����غ�k���9}r�'C�> 3�>�q�
�˙:$�:���9�Ǝ*������m�H�k�����RT.�@��>�F�I*a��1�>s�_��&oԒ������D����ﵳVƏ����<��W���(G�u�v��.b��1 z�3Ȗn<J�aA�j5�l�7%�Ö8���s�Uv��(ΣM��`E�иF�",���������Ǚ5�gj��1������.i�(UĬ(�c���dC|:�.�'ᾯX3y�7N<�U�d�~�sϹ�b������ju7~��������4F�K��`�)}#ֈ���M��C+�<H�H��̨V�?�f��	�x��^.E0:�є7�9�(R����lp�m"��7u]>�#�r����&c����o^�� 릛����߄�g٨�2��R�2�/5'��v��
@-�V*��d��QI�
f�〽c-�rP�kb��&g�n!�H�b̡�4�� ��#�`��3~ uɦ��z�öAH�۰���ߪ��/EPAc��l~O��H�M�V�`�E+5C��ť���x�i>��M G��,\<�F�	���B�7	���_�3���F����$g���K�`/�.rjc���Z�����aO���O^6n&���C��]���M�=maE�NG�����0�*l���g���Fe��;(V��h���?��;ާVny�e�!mW�qRZ|a:�W����{)
*���{ ڃ5*�A�/���ZqS� ��Lj8E0 �S~�h��~�%�#{���x|9����-<?�WH}��^Wf؈%���~и�Xc��L�q>t�*źd �ך�k����Og��_�.�}ֈ�]!�O!�E�����@�F�Z�x)�|�����'��z�b�z������ѿK¹;o㖓Ԟpd��.�JO����o�����s�)Lc��"��֦.�l�C5��P\� ���Pd��tg��nf޹P:sl���O���G؞�D��������͜	���%�������6�wm�t}�����J7̏`�t���֗[3|�JD� ��E�N�ܪ���8�l��\�g}q"�#��f��pP)B��6Kr���=���B��}l}��y�uk≭G? �"OY?DSn����es�j��1_��z�����e�t%�
4�?��h��K\9p�aF+�Hlj��+�Yy/����>� !���:7���=̷a4�7jG��ɭe�zi�Ģ���;���s͞[E�/u%G0/�S�?l!�N�f ^_���w�yW�1}�� |�߷�#�y� ���=��E�Es�_DFS�5�gs����8+��iZn�=�4��Bw�(pM�3]��y�A?�$7�����n�p���VVy��zv��:������h�F�uH�F6r�n99
��N��<�V��	h��Z�a�cx�.
g��h��K& ��MU��S������#k6�"��~}��3!?6R�Am�=f�;hm�t�z�M7��a�O j�3j�ٲ,!G��=�~�,4�+�Fz��M�ȪVP��Z��"�������XZ6%,d@��X�vu�X��� J[!ZB�Cѷ8R˿�M�G|������G/�(���NInr�A�X�턘2دeK �Ǿ�0(� &��*��]P$Rz�`����C����	�)��uV��Q������+F ��a��fC���7-�[��I*s_��G��\﵋����8�H�>�O1��4%{��Zh2uo*��M���t���#E%�7O���C����R뷬��C�>w���rI�J��H2m�xa�m��ÐG��!�לc��	�S�1�O�0#��s/��S���U�-[%��T/L���O"�i7Z�m�к�ŏ*f�gߛĸ3��f�,��Sh����v�d)��յ0��\8�����y��#��΋�������zS�l���;>�i>��z=�u%��c�g�YZ��,�|4�j]���-��L�E�,r�p��Ŵ�q�<	�����qN�jQ`��ť���,}��r�V��F��?�����Y �u������n2�Tֱk������4\���D������5�Ư��]�E�2�R��gc�1T�J���0tyy!���TK3:<�KHخ�P�Ŀbͼ#lW֌�oi������s�Jt�<R�)i*��
�N��>Tk5<'��p�x��j94��8��:Cm�}��5c�D�M�*���7��m�|=�����Q돯ԥLӕ~����w��۴����%�&$�RvU�U.�0�%9~��+&���j��Ղؐ�O����Rh�,I�jc�5�}�Ǽs@��ٛ�]�����%����zUi_�ƅ�H��px5�A��HN��
b�]R���+�"�s�g�
��'��Y4H��4�����'Li�&��\p}"��x�6hv;�1Ox����*�J����g5��!w������ ��&���h��h���S��j�$qLé2����8�Q���2�YrΉ��y��z��$8qY-��.�)j��㉠����5��L�65S�Y���`��6#��?��C`Y*���� �6�����^9�nHR9��J}NoQ]זP�y�,���~qW�"�ľ-]!�?����0�=��~�-
*��A��m�|jk�dtx�����Y�/!ב()�7��m��Zp��&c��@�>�����S�x�ք�g��oHܜ�����1�+Yi���w��xk󲍾�󗂺p{I-�e�/��֛�
�p(�z9�����W6&U` �^���iIx�r�oZ�D�ӠU%w�)����*x��p��X�o�RD&�*�zD��3���Y��G;�#K�8��N
p�������5�՛�/Ȯ�w���;-�Pp�_���
bXZ���G̵U1��)a�N�:;D�t���UC)���/�g��Q�ӌZ����^ږ�@M#��{�P����y�<���W�w��������� ����V�y$�n���`.nU�8L���k���s���{��mG}�VW.�5_o ��ڵ�̔��a��˾6���S��"!�Hk�Zm_"��3_}.N���Z��1�����u���c�p�z����	u��o�6��!���$���b��L�lJDǆ����c���~����P��wN��H��IT9/��-d�S��L���AP4g�Q�y͕�^�9����3� a�:??�B?J
�[a���Mp>Q.h���L_��X����.w��o�[Ơ��Q�g;��2�
c�O!nC?��x���4����m�����c�r����J8z����iJ4�F�������1+I܏&����M"���ҧ�?;UO�SXlxVHYEB    4f62     b50
HAv��=0��g`�B�'�=�4� h��_���L&v����nܳ���C�wo����]�t���9����i�F"����:;�V��T�M�t��o
�볹�^�	�7�#;c�bJ ������p���tb�|r���C�npx��)�?�����3���v7��bIH�E��e]TGwdb�˶M��v@3�����P��-�q����$�'4�e2�Buwe�~��KQs<k����#����9����nh������#�p�4��~;J�*��Spk�w. ���,��#OO�A���?����/9j��g���WG��fK""&�@�s�oٴ���e��;�X��"k��ke4�g�X���[	r��5:U�U�����T׮1I�酼"�ٳ���:�;�4L��N�*,eW<�lqq<(�M#+����Kʵ�]g�^���
xayե�fU3���ኈ�J�@wsz^Qʌ�X&���n!v"F�D���$]�6���H��h$�<�3�Q�QV:�i�A_�#���?�nD};q�����-�<�
�)�=�ƞ��[��$%]�?�q���fn髌���x><%�tx��oO��V(����O�����|ظO\=��o2�Տ#�$`ΐ���!��0��Ϫs�XY� 7�%j񐱄�����NnU����a���w]H�n�R�ܝ݈6�$O�'c�:���&��.���H!*~�'����,�V��;��8 �蚔��B��7`�K�X�����ۙ��]�Fl�E��V��h��υJYN=t�[֧w����@��f�v����j
':lױ���u,4~aPhV���P���F3b	����ϣ곖 �t�Ԭ���E�lJ-G�w�á4�7�A���3WM� #gr�^���K�v!�������`F�� d)E#��
_86�nr�I
ıR�}õ� ���3�)��;�q�O���
����E�9�����ԅ��P�б~x�`���<��cf�5��y�j�0%v9��G��
��:𛔝ΐg���ȼ4�M �qI	6��q�� Y.���J�qh�e�R(��unAOS�lۀe��cy�A}*i+ΒL��@����t��
��˳�*l&�gK�����O�
TzsO	.ㇹ�.2��h�TY�HhƷϷJvi*9��w���Mݲ��HK�k�d�/װ:U�	L���)�*���%��a�r}i5�h��L���׎���0�+��i�T�;��3��>G�`P�3�VI,;�������s��(-,i��3��uD�M�i�"��L��T�u�8gO���~�q(L�*c�/��b"
4��B�ck�Z�(b��?�jwm�������@k�[n��������]g�Wdu|���x��mi'�P��r�r����V���a��;�dS&��,��7�j�dr�E�i@�iRQo��? �h
]�Y"⹿�%E��
���l^�Q�Ҁ8�	i��Mw'8�`څ�D���h 	r �^V�{���&�8�@Sw
����o�F�nr�L��Tv�MMԝ���ȎH�i���ќ�Z�xs�T���˘����~�<%��= щV����G4j{)F_9;�`7�jv�'q�m��k��+���}��-j�N��w�`|�M�{}	���z�0���E:J�ڇ�{�E��Ǆ�fM0�i�4���qs}"8Ro%�5�.��*���H�kg���V�/TX���7]b���fKs�W�ř^�A9���.���Z3�~V2�~�Nb�s �����ܢ?�aEvE�ŴR^���T��@g.S"˙�:m�W�ur ��s(��2����GP#U+��͆w��'ջ�������'W�م��a�^_���(����໗H�=��g�(Z�t���6:w�3 k�zuSBcgl<�0�~}8mj�S��`i�
8�fZ�X>�%k�I	[�t���I�G��2|��z| &�౫ΗA&�;'�4f��!�Q|GX!�&j�R��=�^,����3�k)�Ê�bTic�Ca�oM�Ε=-���x�l��&���uQ队���BS�3�*H�u��W^n�g.Ґj�z�(PB���2��(����ƩX�e��3ڙz��$�,ZQPv�!u���y�Z�$���9��]�yW�Ů✰��5ڳ,����lGW7��?�ZE�S,e��D�F<zdS_�`�Cf\��$�h�&�*�5NcY�A�٢�_z?q|ٚ>頺F��J�K�j���#ϕ���8m�n�7�e�6kY��f@��
y���ɲ�56y9�Ϩ��pa�h��nH]Qq��cx�[N�q��j����G!Z{����n�܎X����R�]�S��$�3ʉr���^x�ﰬ�f���� ��Ѐ���=�1��
�g�a@e2��)x5����_�6^".�?��XW�|����e.f�.%������UM�	o�}�%�g��>�ѿa��)�8&NJ*��w=��u��l���?� [}��7^��h.�=6�pp�J ��D�zA����y��r�­\(�g�����n$h�ic;�q����c*:�S�N媍R|�i16��2������ke��8=
�	��$�Jw|Z�ĵ֦��jw��Ÿ��_��$/�����-��D��J��  i9��"o+�]���0^�^��~��a]�/"��*�\���5�A����-lx�4��<@���r�O�j����Pw1I��/&�W����E"]����M�R#߬�Z2	���Y�k�{S^B�,�3�Sp^=�y����8F;�-Gӊ���}F�2�<׳Z"!vT:�����iq� @��Rh5���9�㫽<�8'��ύ:*7e�