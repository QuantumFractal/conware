XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���:IIo9��
I���L��s�T�H���6,��%q�~R��!��Q�,\l�V�Z��	�`�0�Z���み~&�i���+P�A��	��
o�B���g���7,4�b��HḀb�q���|���޶��4����L�Z9��{e��\�����PM@�߆�2,����I�uV�]�*��q؇��Em��r�ȋ1r�O�@�8Ph:����Th
�i0����ɕ�Bk���Du�"{hs��rX����U��%ҏN�J�R��̱ϒ�2��h<)�hYc�����"�R}Gϰ\J�$��[(����2�Z��C&�i�B�V��Tﲝ�'2l`���#�2���{�:3�Z1��b���y�ω[�@O�n"��߬]I���/�j����@Qǃd}������[��0��ߊ1<�# 9636U���OsGԥ泎����Z�0L�sb�[�������Fh��9��벪�_��@�ԩ�m�վ��d�<�2N��^��:t��&���r�c��!J�ȭ�W���@ž� /�ͦ�h�"�/��'z���$�U���ϛ߶� ?�%�ֵɮ�L�q�$�l����b�ߊWn_���Դa�h��~�ϱ�s�lxo�UN�r�}^�g�#Q:�g����Z�f$�-�uO�|LfIMK��Q�E�h�.�j���'��Q�H���HT��t/�����4{�v��}_&����z��{U'���h�I�uD�����u|<�������}r�XlxVHYEB     f6d     6f0E�}��8�L�$4`Z��ʽ�+��Y��J���a��@�����-9�s��:�<�5"_�I�X���TR�����Dﶶ�<�'�����.��8���Pw��xG2zT|#�ջ����\z�v�����h�mv�v��2����E<ߔ�
	}��w����D@��T�6{D���R�]{�gQ
�̖9 ������+̭��2e8&��3eu�:Nɷ�}��8�JZrԒ�2 ܑ�z�_=��_�6����+��K���d8��z�E��x��e�[b�
/�,����S�����+���I�RU@��G�sP�+Z%��\�#��O�y���+���[��筓r�'���7��$����;�@�q4c�:��`a�n���Еp�GsyI1���!|���a2�&_�|�����;��?�����&�q�7/R1��Tm�6g��M�E�2�pG�3鷕X����L�v�&���6m�΍��?҃�9�>���W���%@�լ�L��A{W��}�TF����hC�
�X�{��_XV�·��R-��3�2�|}�c.��F�)� �<�j���_~�G�& ��#h �f�b�)=�mD���s��r��? J/�)�)����η����9�z�>?r2�ٚ���eDS3��'��-�
�^��+�eaY��xT��[���E��>�%E��<������x�'��������#�l �(�~�L$���{��|86#젅��8X������گq4���P�f2���=6��,/G.���BU6�om�)��VQ��÷U��m0�ՈyV����"���u,U2m��$k�Vl��3�w��"*�G���,�f2OG�־�+V�v����g�;�q�dˈ�o�����byF��R��iL���Tu�d���[:F*��SɃ�^
Q&L-��㦣�	�;� Q���jJ�@�rfGft��z��V�ن�8�;t']��*�w䐘�$�Z�:�zP��qI�#r��*a5�u�<]Hp��9�3�"4��,�Ü2>�����cbw�gg�Q_!�B��<w�5��7�FQ=K#j{��z��+���.Q�> ��Y(�]X���'n���`3����\�D9�E*�)\t4���c2�E�nE�e���kfx�t�G�׋�~���dO1������	���moz�u�2�d�f m"Qg�{E$�.&�05=��霅f�W�#�n;��g�é&3`z�ꨲK���m�e�๥�m�{a�K���}d��K�p����m����	!zg �˧TPڀ��kW��CM�'��o�s�zr�s#��c�g*e�]��7T�h�:� m�O��]j���>Am=F�,Z��ܰ�s��nNW&�0�YD�������������rLD��E�s��ѝv����.ȫ0T�0SZ<Gҭj_K[O���o'Q��wS�U�?Xz!v(7�ELVMtRzo;ܖ�4 R7 ��[�9+]N@��\\,I��F����2RjV���,�臲۱XT��z�K�$��X���'����.=�`���XݬP�lW�ňV�'�"n�ϔ\��[�
��e�a�O�
6�·��~����[��@�9�zu�� N��61#�jf=�hU����qeL����)bi)�x��y�����dF��ܬ6�]���sl����,��2W\��~?{6L��,�����U���z>��rm�C�̓��<tFc��N�T��%y�#�u+c���wÈq\⸜���s�}6���wC�