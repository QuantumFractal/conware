XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��-p^�>��.�6�Y�9�����£؆	M ��IBp��@�`sÔ���V���k�Y���_�6���[p/|�\Q��'�${�;��d)�	�ֲ��I�\)U�?�Ts��BĄ��Tn7�C�q0�y~OU.e>�4C|� ���]�;����#7��h&$C��B%T^	�A����u��1t��/y�b��k �.��=E&v�
V����;��2j�1�/��QeZ�!^]��I!�J�t��Y��>�I�Ǿ��4��ܚ�9�0��q�/��8�x������.���+�r� �������:rH�*�i�첇m�9+0�h�u�z6�}'yk:���Rd�r�( o�%�N�L{M�1�Pa��Y9�
��{�%-jծF�S�܈Ҹ�B�u ��8�HY�:'�zX���8.'E��i���Ƅg�,���}�;���F���`��i��px��^M+�	��"����?�B�T�{�]a+���KM�ŧ��o�8�PV2�_Ζ�Ki%Y����}Y�ꈒ'`���?�9�G,�RK�엔?����Gip�u���?e҉(cW�-�������mYZ3����T~�ھ�z@��gpG^�FkEr*�e����P���h���<����O������e!��H���W8�2���[<�ϱP��.�.�{�Su�|��	����Xq|��:)�"��4�����XH����nN�����j��Q�h�7iʛo�ľf_�rYk�aa4ZO`p�W���7p��E��XlxVHYEB    1853     810�C1�L i����2gtf@����^O.�)�͸���/7K��	F`M�'R(CBߎ��2/�O�O�C�O a4�),�#**3!������w�DLw�M�O�#���c��SU҄nn.��>ܮ#JY�	�~��uL��6�hsu����;��8��~��,O��Ճ'\�F��L����Z�r ?_l'��=5t����"V�R��J����d(+#a�I�[����� ��������<�(�����w��V/e�1�����_0-�|�jK)5;\N{C�*(�/6܇n%��sp�dP��l��p�T���UA�hcl�[<�1���� �C�I�]'�e[��Ώ{3B?�R�6=5�� 7�i(� ,�� *I�D�ʯ�Y�}��0e����1�تȖB$��Ǘ8�H�!�5| ��<�ſ@�u�d$P��<��(�����;���C�̿�|>�hj5�0�	��"�B�,�䑿S���n:m���"�9l��ŝ_QS0/��@6��y����k^��-mp�U)��i�kX�x)�H�?%��Ӷr�u��h�kv�}�����^�Cjm��g2�] ��gq�)�AR6�M��w�V9�� Z����p�V� �8L�$8��Fj��=t�7A��:��c�X��ɱ�v/��ef
�''��;К���j�/�d�b�=��Y��JCw{��7) d�%183��%"-���ٌ1q aPrs\ePO��MRU����m͵�D��⽿�#mkζ�]�e�Q�\�ۯ�j+�-��S��i]�.20�z&|��\1< C��e�,���Dz���BQ��u��G��9
 �-�;:�ޮ���	5�i�0��t��1�H&�fR`y�
.?6YY%�$+7*�As�q:4�N�vf���R����po�ny��_�pda�,L�Bu^b�?�e�U>�zm�ͣ��M�&�Ð|IB��G���j6:�,-��t�봪o�j&&�����	Kb�Г]L3�!��!�ݥ�)�<7���I�QQm�>���L�2n�E�H>I�>���)���;n���:0j��
)�0�ƸdϠ-��ܡOf��u�߄
I�5Z@�TTh�yLxn�I��[Dk���������������d|�,i�W֊U�NM}�Ŀ�^(�ġ������if��`�D�ݍ��Y�`l(in�q�����vS�:�z����p	�	K��@0��z�E��_�����]�=l]&ɌW�;NP��������ѬҴ'��i�ܿ����UiCþٷ#����#/�l�%p<l��e�?�L55-���P��Ȅ��و���+�p5�a��D��zn��8$�3�]�T��9X-��̰L�Ԥ+Ri뺉���
(�_*t0��[bd~`)����3ߨ<�N4���:�O9��iz_})����y7��p;nl'�e7Ӿ�:dg��뙷-WhF�Zó_t�;^6F�9�nA�N���v�:�~%��j��KhاRc!eB����s�n�g����1�����&��ɸ��jE�@.��2��l��g-�@|��J3��Ŀ3Sp)�վ&T����ka-�FL�+W�|�A4-qWQ�[����*dX^3��d����=�Po��m����e;�|�(��Z�j&E|�lJ~��P�`��k5�Q ¶����e��Ć���:*�B�|�vX��Aꒀ9�6� 5��^�C�F�<�D���V����ǻ� ��aj��M/���x�H���jTC��9��9)�*��w�D�T�6c�)xҹ	� ���pK�K�J�BؽC��_9��`H"[K�����hj�MI����/�M�KW�K�o�s�K^a!F�a�nm�r�@�:*��EK�(r�ki�|�n 
$@&�}br��\�o���;�H\! ��:��8��P�9����1 �k��}�,P-��`y\���W;�R�\Q~u�"#�N����*2�h��؅ ���%���T�R;/�T:`�T(�-���i�.�OU�
p�@ɏ޳�N